//------------------------------------------------------------------------------
// The confidential and proprietary information contained in this file may
// only be used by a person authorised under and to the extent permitted
// by a subsisting licensing agreement from ARM Limited.
//
//            (C) COPYRIGHT 2010-2015 ARM Limited.
//                ALL RIGHTS RESERVED
//
// This entire notice must be reproduced on all copies of this file
// and copies of this file may only be made by a person if such person is
// permitted to do so under the terms of a subsisting license agreement
// from ARM Limited.
//
//      SVN Information
//
//      Checked In          : $Date: 2015-09-22 12:44:46 +0100 (Tue, 22 Sep 2015) $
//
//      Revision            : $Revision: 320568 $
//
//      Release Information : Cortex-M0 DesignStart-r1p0-00rel0
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Cortex-M0 DesignStart processor logic level
//------------------------------------------------------------------------------

module cortexm0ds_logic
(hclk, hreset_n, haddr_o, hburst_o, hmastlock_o, hprot_o,
hsize_o, htrans_o, hwdata_o, hwrite_o, hrdata_i, hready_i, hresp_i,
nmi_i, irq_i, txev_o, rxev_i, lockup_o, sys_reset_req_o, st_clk_en_i,
st_calib_i, sleeping_o, vis_r0_o, vis_r1_o, vis_r2_o, vis_r3_o, vis_r4_o
, vis_r5_o, vis_r6_o, vis_r7_o, vis_r8_o, vis_r9_o, vis_r10_o, vis_r11_o
, vis_r12_o, vis_r14_o, vis_msp_o, vis_psp_o, vis_pc_o, vis_apsr_o,
vis_tbit_o, vis_ipsr_o, vis_control_o, vis_primask_o);

output [31:0] haddr_o;
output [2:0] hburst_o;
output [3:0] hprot_o;
output [2:0] hsize_o;
output [1:0] htrans_o;
output [31:0] hwdata_o;
input [31:0] hrdata_i;
input [31:0] irq_i;
input [25:0] st_calib_i;
output [31:0] vis_r0_o;
output [31:0] vis_r1_o;
output [31:0] vis_r2_o;
output [31:0] vis_r3_o;
output [31:0] vis_r4_o;
output [31:0] vis_r5_o;
output [31:0] vis_r6_o;
output [31:0] vis_r7_o;
output [31:0] vis_r8_o;
output [31:0] vis_r9_o;
output [31:0] vis_r10_o;
output [31:0] vis_r11_o;
output [31:0] vis_r12_o;
output [31:0] vis_r14_o;
output [29:0] vis_msp_o;
output [29:0] vis_psp_o;
output [30:0] vis_pc_o;
output [3:0] vis_apsr_o;
output [5:0] vis_ipsr_o;
input hclk;
input hreset_n;
input hready_i;
input hresp_i;
input nmi_i;
input rxev_i;
input st_clk_en_i;
output hmastlock_o;
output hwrite_o;
output txev_o;
output lockup_o;
output sys_reset_req_o;
output sleeping_o;
output vis_tbit_o;
output vis_control_o;
output vis_primask_o;

wire Lnh675, Doh675, Hph675, Jqh675, Lrh675, Lsh675, Tth675, Bvh675, Gwh675, Oxh675;
wire Wyh675, E0i675, M1i675, U2i675, C4i675, G5i675, N6i675, T7i675, A9i675, Hai675;
wire Obi675, Vci675, Cei675, Jfi675, Qgi675, Xhi675, Eji675, Lki675, Tli675, Bni675;
wire Joi675, Rpi675, Zqi675, Hsi675, Lti675, Pui675, Tvi675, Xwi675, Byi675, Fzi675;
wire J0j675, N1j675, R2j675, V3j675, A5j675, F6j675, I7j675, L8j675, O9j675, Raj675;
wire Ubj675, Xcj675, Aej675, Dfj675, Ggj675, Jhj675, Mij675, Pjj675, Skj675, Vlj675;
wire Ymj675, Boj675, Epj675, Hqj675, Krj675, Nsj675, Qtj675, Tuj675, Wvj675, Zwj675;
wire Cyj675, Fzj675, I0k675, K1k675, M2k675, O3k675, Q4k675, S5k675, U6k675, W7k675;
wire D9k675, Nak675, Ybk675, Idk675, Sek675, Cgk675, Mhk675, Wik675, Gkk675, Qlk675;
wire Ank675, Kok675, Upk675, Frk675, Qsk675, Buk675, Mvk675, Xwk675, Iyk675, Tzk675;
wire E1l675, P2l675, A4l675, L5l675, W6l675, H8l675, S9l675, Dbl675, Ocl675, Zdl675;
wire Kfl675, Vgl675, Gil675, Rjl675, Cll675, Mml675, Wnl675, Gpl675, Qql675, Asl675;
wire Ktl675, Uul675, Ewl675, Oxl675, Yyl675, J0m675, U1m675, F3m675, Q4m675, B6m675;
wire M7m675, X8m675, Iam675, Tbm675, Edm675, Pem675, Agm675, Lhm675, Wim675, Hkm675;
wire Slm675, Dnm675, Oom675, Zpm675, Krm675, Vsm675, Gum675, Nvm675, Xwm675, Jym675;
wire Vzm675, H1n675, T2n675, F4n675, R5n675, D7n675, P8n675, Z9n675, Jbn675, Tcn675;
wire Den675, Nfn675, Xgn675, Hin675, Rjn675, Bln675, Lmn675, Vnn675, Gpn675, Rqn675;
wire Csn675, Ntn675, Yun675, Jwn675, Uxn675, Ezn675, O0o675, Y1o675, I3o675, S4o675;
wire C6o675, M7o675, W8o675, Gao675, Qbo675, Bdo675, Meo675, Xfo675, Iho675, Tio675;
wire Eko675, Plo675, Zmo675, Hoo675, Spo675, Aro675, Iso675, Rto675, Gvo675, Mwo675;
wire Vxo675, Ezo675, N0p675, W1p675, F3p675, O4p675, X5p675, J7p675, V8p675, Fap675;
wire Nbp675, Wcp675, Cep675, Ifp675, Ogp675, Uhp675, Gjp675, Skp675, Amp675, Pnp675;
wire Epp675, Tqp675, Isp675, Xtp675, Mvp675, Bxp675, Qyp675, F0q675, U1q675, K3q675;
wire A5q675, Q6q675, G8q675, W9q675, Mbq675, Cdq675, Seq675, Igq675, Yhq675, Ojq675;
wire Elq675, Umq675, Koq675, Aqq675, Qrq675, Gtq675, Wuq675, Mwq675, Cyq675, Szq675;
wire I1r675, S2r675, F4r675, S5r675, E7r675, O8r675, Aar675, Mbr675, Ycr675, Ker675;
wire Wfr675, Dgr675, Kgr675, Rgr675, Ygr675, Fhr675, Mhr675, Thr675, Air675, Hir675;
wire Oir675, Vir675, Cjr675, Jjr675, Qjr675, Xjr675, Ekr675, Lkr675, Skr675, Zkr675;
wire Glr675, Nlr675, Ulr675, Bmr675, Imr675, Pmr675, Wmr675, Dnr675, Knr675, Rnr675;
wire Ynr675, For675, Mor675, Tor675, Apr675, Hpr675, Opr675, Vpr675, Cqr675, Jqr675;
wire Qqr675, Xqr675, Err675, Lrr675, Srr675, Zrr675, Gsr675, Nsr675, Usr675, Btr675;
wire Itr675, Ptr675, Wtr675, Dur675, Kur675, Rur675, Yur675, Fvr675, Mvr675, Tvr675;
wire Awr675, Hwr675, Owr675, Vwr675, Cxr675, Jxr675, Qxr675, Xxr675, Eyr675, Lyr675;
wire Syr675, Zyr675, Gzr675, Nzr675, Uzr675, B0s675, I0s675, P0s675, W0s675, D1s675;
wire K1s675, R1s675, Y1s675, F2s675, M2s675, T2s675, A3s675, H3s675, O3s675, V3s675;
wire C4s675, J4s675, Q4s675, X4s675, E5s675, L5s675, S5s675, Z5s675, G6s675, N6s675;
wire U6s675, B7s675, I7s675, P7s675, W7s675, D8s675, K8s675, R8s675, Y8s675, F9s675;
wire M9s675, T9s675, Aas675, Has675, Oas675, Vas675, Cbs675, Jbs675, Qbs675, Xbs675;
wire Ecs675, Lcs675, Scs675, Zcs675, Gds675, Nds675, Uds675, Bes675, Ies675, Pes675;
wire Wes675, Dfs675, Kfs675, Rfs675, Yfs675, Fgs675, Mgs675, Tgs675, Ahs675, Hhs675;
wire Ohs675, Vhs675, Cis675, Jis675, Qis675, Xis675, Ejs675, Ljs675, Sjs675, Zjs675;
wire Gks675, Nks675, Uks675, Bls675, Ils675, Pls675, Wls675, Dms675, Kms675, Rms675;
wire Yms675, Fns675, Mns675, Tns675, Aos675, Hos675, Oos675, Vos675, Cps675, Jps675;
wire Qps675, Xps675, Eqs675, Lqs675, Sqs675, Zqs675, Grs675, Nrs675, Urs675, Bss675;
wire Iss675, Pss675, Wss675, Dts675, Kts675, Rts675, Yts675, Fus675, Mus675, Tus675;
wire Avs675, Hvs675, Ovs675, Vvs675, Cws675, Jws675, Qws675, Xws675, Exs675, Lxs675;
wire Sxs675, Zxs675, Gys675, Nys675, Uys675, Bzs675, Izs675, Pzs675, Wzs675, D0t675;
wire K0t675, R0t675, Y0t675, F1t675, M1t675, T1t675, A2t675, H2t675, O2t675, V2t675;
wire C3t675, J3t675, Q3t675, X3t675, E4t675, L4t675, S4t675, Z4t675, G5t675, N5t675;
wire U5t675, B6t675, I6t675, P6t675, W6t675, D7t675, K7t675, R7t675, Y7t675, F8t675;
wire M8t675, T8t675, A9t675, H9t675, O9t675, V9t675, Cat675, Jat675, Qat675, Xat675;
wire Ebt675, Lbt675, Sbt675, Zbt675, Gct675, Nct675, Uct675, Bdt675, Idt675, Pdt675;
wire Wdt675, Det675, Ket675, Ret675, Yet675, Fft675, Mft675, Tft675, Agt675, Hgt675;
wire Ogt675, Vgt675, Cht675, Jht675, Qht675, Xht675, Eit675, Lit675, Sit675, Zit675;
wire Gjt675, Njt675, Ujt675, Bkt675, Ikt675, Pkt675, Wkt675, Dlt675, Klt675, Rlt675;
wire Ylt675, Fmt675, Mmt675, Tmt675, Ant675, Hnt675, Ont675, Vnt675, Cot675, Jot675;
wire Qot675, Xot675, Ept675, Lpt675, Spt675, Zpt675, Gqt675, Nqt675, Uqt675, Brt675;
wire Irt675, Prt675, Wrt675, Dst675, Kst675, Rst675, Yst675, Ftt675, Mtt675, Ttt675;
wire Aut675, Hut675, Out675, Vut675, Cvt675, Jvt675, Qvt675, Xvt675, Ewt675, Lwt675;
wire Swt675, Zwt675, Gxt675, Nxt675, Uxt675, Byt675, Iyt675, Pyt675, Wyt675, Dzt675;
wire Kzt675, Rzt675, Yzt675, F0u675, M0u675, T0u675, A1u675, H1u675, O1u675, V1u675;
wire C2u675, J2u675, Q2u675, X2u675, E3u675, L3u675, S3u675, Z3u675, G4u675, N4u675;
wire U4u675, B5u675, I5u675, P5u675, W5u675, D6u675, K6u675, R6u675, Y6u675, F7u675;
wire M7u675, T7u675, A8u675, H8u675, O8u675, V8u675, C9u675, J9u675, Q9u675, X9u675;
wire Eau675, Lau675, Sau675, Zau675, Gbu675, Nbu675, Ubu675, Bcu675, Icu675, Pcu675;
wire Wcu675, Ddu675, Kdu675, Rdu675, Ydu675, Feu675, Meu675, Teu675, Afu675, Hfu675;
wire Ofu675, Vfu675, Cgu675, Jgu675, Qgu675, Xgu675, Ehu675, Lhu675, Shu675, Zhu675;
wire Giu675, Niu675, Uiu675, Bju675, Iju675, Pju675, Wju675, Dku675, Kku675, Rku675;
wire Yku675, Flu675, Mlu675, Tlu675, Amu675, Hmu675, Omu675, Vmu675, Cnu675, Jnu675;
wire Qnu675, Xnu675, Eou675, Lou675, Sou675, Zou675, Gpu675, Npu675, Upu675, Bqu675;
wire Iqu675, Pqu675, Wqu675, Dru675, Kru675, Rru675, Yru675, Fsu675, Msu675, Tsu675;
wire Atu675, Htu675, Otu675, Vtu675, Cuu675, Juu675, Quu675, Xuu675, Evu675, Lvu675;
wire Svu675, Zvu675, Gwu675, Nwu675, Uwu675, Bxu675, Ixu675, Pxu675, Wxu675, Dyu675;
wire Kyu675, Ryu675, Yyu675, Fzu675, Mzu675, Tzu675, A0v675, H0v675, O0v675, V0v675;
wire C1v675, J1v675, Q1v675, X1v675, E2v675, L2v675, S2v675, Z2v675, G3v675, N3v675;
wire U3v675, B4v675, I4v675, P4v675, W4v675, D5v675, K5v675, R5v675, Y5v675, F6v675;
wire M6v675, T6v675, A7v675, H7v675, O7v675, V7v675, C8v675, J8v675, Q8v675, X8v675;
wire E9v675, L9v675, S9v675, Z9v675, Gav675, Nav675, Uav675, Bbv675, Ibv675, Pbv675;
wire Wbv675, Dcv675, Kcv675, Rcv675, Ycv675, Fdv675, Mdv675, Tdv675, Aev675, Hev675;
wire Oev675, Vev675, Cfv675, Jfv675, Qfv675, Xfv675, Egv675, Lgv675, Sgv675, Zgv675;
wire Ghv675, Nhv675, Uhv675, Biv675, Iiv675, Piv675, Wiv675, Djv675, Kjv675, Rjv675;
wire Yjv675, Fkv675, Mkv675, Tkv675, Alv675, Hlv675, Olv675, Vlv675, Cmv675, Jmv675;
wire Qmv675, Xmv675, Env675, Lnv675, Snv675, Znv675, Gov675, Nov675, Uov675, Bpv675;
wire Ipv675, Ppv675, Wpv675, Dqv675, Kqv675, Rqv675, Yqv675, Frv675, Mrv675, Trv675;
wire Asv675, Hsv675, Osv675, Vsv675, Ctv675, Jtv675, Qtv675, Xtv675, Euv675, Luv675;
wire Suv675, Zuv675, Gvv675, Nvv675, Uvv675, Bwv675, Iwv675, Pwv675, Wwv675, Dxv675;
wire Kxv675, Rxv675, Yxv675, Fyv675, Myv675, Tyv675, Azv675, Hzv675, Ozv675, Vzv675;
wire C0w675, J0w675, Q0w675, X0w675, E1w675, L1w675, S1w675, Z1w675, G2w675, N2w675;
wire U2w675, B3w675, I3w675, P3w675, W3w675, D4w675, K4w675, R4w675, Y4w675, F5w675;
wire M5w675, T5w675, A6w675, H6w675, O6w675, V6w675, C7w675, J7w675, Q7w675, X7w675;
wire E8w675, L8w675, S8w675, Z8w675, G9w675, N9w675, U9w675, Baw675, Iaw675, Paw675;
wire Waw675, Dbw675, Kbw675, Rbw675, Ybw675, Fcw675, Mcw675, Tcw675, Adw675, Hdw675;
wire Odw675, Vdw675, Cew675, Jew675, Qew675, Xew675, Efw675, Lfw675, Sfw675, Zfw675;
wire Ggw675, Ngw675, Ugw675, Bhw675, Ihw675, Phw675, Whw675, Diw675, Kiw675, Riw675;
wire Yiw675, Fjw675, Mjw675, Tjw675, Akw675, Hkw675, Okw675, Vkw675, Clw675, Jlw675;
wire Qlw675, Xlw675, Emw675, Lmw675, Smw675, Zmw675, Gnw675, Nnw675, Unw675, Bow675;
wire Iow675, Pow675, Wow675, Dpw675, Kpw675, Rpw675, Ypw675, Fqw675, Mqw675, Tqw675;
wire Arw675, Hrw675, Orw675, Vrw675, Csw675, Jsw675, Qsw675, Xsw675, Etw675, Ltw675;
wire Stw675, Ztw675, Guw675, Nuw675, Uuw675, Bvw675, Ivw675, Pvw675, Wvw675, Dww675;
wire Kww675, Rww675, Yww675, Fxw675, Mxw675, Txw675, Ayw675, Hyw675, Oyw675, Vyw675;
wire Czw675, Jzw675, Qzw675, Xzw675, E0x675, L0x675, S0x675, Z0x675, G1x675, N1x675;
wire U1x675, B2x675, I2x675, P2x675, W2x675, D3x675, K3x675, R3x675, Y3x675, F4x675;
wire M4x675, T4x675, A5x675, H5x675, O5x675, V5x675, C6x675, J6x675, Q6x675, X6x675;
wire E7x675, L7x675, S7x675, Z7x675, G8x675, N8x675, U8x675, B9x675, I9x675, P9x675;
wire W9x675, Dax675, Kax675, Rax675, Yax675, Fbx675, Mbx675, Tbx675, Acx675, Hcx675;
wire Ocx675, Vcx675, Cdx675, Jdx675, Qdx675, Xdx675, Eex675, Lex675, Sex675, Zex675;
wire Gfx675, Nfx675, Ufx675, Bgx675, Igx675, Pgx675, Wgx675, Dhx675, Khx675, Rhx675;
wire Yhx675, Fix675, Mix675, Tix675, Ajx675, Hjx675, Ojx675, Vjx675, Ckx675, Jkx675;
wire Qkx675, Xkx675, Elx675, Llx675, Slx675, Zlx675, Gmx675, Nmx675, Umx675, Bnx675;
wire Inx675, Pnx675, Wnx675, Dox675, Kox675, Rox675, Yox675, Fpx675, Mpx675, Tpx675;
wire Aqx675, Hqx675, Oqx675, Vqx675, Crx675, Jrx675, Qrx675, Xrx675, Esx675, Lsx675;
wire Ssx675, Zsx675, Gtx675, Ntx675, Utx675, Bux675, Iux675, Pux675, Wux675, Dvx675;
wire Kvx675, Rvx675, Yvx675, Fwx675, Mwx675, Twx675, Axx675, Hxx675, Oxx675, Vxx675;
wire Cyx675, Jyx675, Qyx675, Xyx675, Ezx675, Lzx675, Szx675, Zzx675, G0y675, N0y675;
wire U0y675, B1y675, I1y675, P1y675, W1y675, D2y675, K2y675, R2y675, Y2y675, F3y675;
wire M3y675, T3y675, A4y675, H4y675, O4y675, V4y675, C5y675, J5y675, Q5y675, X5y675;
wire E6y675, L6y675, S6y675, Z6y675, G7y675, N7y675, U7y675, B8y675, I8y675, P8y675;
wire W8y675, D9y675, K9y675, R9y675, Y9y675, Fay675, May675, Tay675, Aby675, Hby675;
wire Oby675, Vby675, Ccy675, Jcy675, Qcy675, Xcy675, Edy675, Ldy675, Sdy675, Zdy675;
wire Gey675, Ney675, Uey675, Bfy675, Ify675, Pfy675, Wfy675, Dgy675, Kgy675, Rgy675;
wire Ygy675, Fhy675, Mhy675, Thy675, Aiy675, Hiy675, Oiy675, Viy675, Cjy675, Jjy675;
wire Qjy675, Xjy675, Eky675, Lky675, Sky675, Zky675, Gly675, Nly675, Uly675, Bmy675;
wire Imy675, Pmy675, Wmy675, Dny675, Kny675, Rny675, Yny675, Foy675, Moy675, Toy675;
wire Apy675, Hpy675, Opy675, Vpy675, Cqy675, Jqy675, Qqy675, Xqy675, Ery675, Lry675;
wire Sry675, Zry675, Gsy675, Nsy675, Usy675, Bty675, Ity675, Pty675, Wty675, Duy675;
wire Kuy675, Ruy675, Yuy675, Fvy675, Mvy675, Tvy675, Awy675, Hwy675, Owy675, Vwy675;
wire Cxy675, Jxy675, Qxy675, Xxy675, Eyy675, Lyy675, Syy675, Zyy675, Gzy675, Nzy675;
wire Uzy675, B0z675, I0z675, P0z675, W0z675, D1z675, K1z675, R1z675, Y1z675, F2z675;
wire M2z675, T2z675, A3z675, H3z675, O3z675, V3z675, C4z675, J4z675, Q4z675, X4z675;
wire E5z675, L5z675, S5z675, Z5z675, G6z675, N6z675, U6z675, B7z675, I7z675, P7z675;
wire W7z675, D8z675, K8z675, R8z675, Y8z675, F9z675, M9z675, T9z675, Aaz675, Haz675;
wire Oaz675, Vaz675, Cbz675, Jbz675, Qbz675, Xbz675, Ecz675, Lcz675, Scz675, Zcz675;
wire Gdz675, Ndz675, Udz675, Bez675, Iez675, Pez675, Wez675, Dfz675, Kfz675, Rfz675;
wire Yfz675, Fgz675, Mgz675, Tgz675, Ahz675, Hhz675, Ohz675, Vhz675, Ciz675, Jiz675;
wire Qiz675, Xiz675, Ejz675, Ljz675, Sjz675, Zjz675, Gkz675, Nkz675, Ukz675, Blz675;
wire Ilz675, Plz675, Wlz675, Dmz675, Kmz675, Rmz675, Ymz675, Fnz675, Mnz675, Tnz675;
wire Aoz675, Hoz675, Ooz675, Voz675, Cpz675, Jpz675, Qpz675, Xpz675, Eqz675, Lqz675;
wire Sqz675, Zqz675, Grz675, Nrz675, Urz675, Bsz675, Isz675, Psz675, Wsz675, Dtz675;
wire Ktz675, Rtz675, Ytz675, Fuz675, Muz675, Tuz675, Avz675, Hvz675, Ovz675, Vvz675;
wire Cwz675, Jwz675, Qwz675, Xwz675, Exz675, Lxz675, Sxz675, Zxz675, Gyz675, Nyz675;
wire Uyz675, Bzz675, Izz675, Pzz675, Wzz675, D00775, K00775, R00775, Y00775, F10775;
wire M10775, T10775, A20775, H20775, O20775, V20775, C30775, J30775, Q30775, X30775;
wire E40775, L40775, S40775, Z40775, G50775, N50775, U50775, B60775, I60775, P60775;
wire W60775, D70775, K70775, R70775, Y70775, F80775, M80775, T80775, A90775, H90775;
wire O90775, V90775, Ca0775, Ja0775, Qa0775, Xa0775, Eb0775, Lb0775, Sb0775, Zb0775;
wire Gc0775, Nc0775, Uc0775, Bd0775, Id0775, Pd0775, Wd0775, De0775, Ke0775, Re0775;
wire Ye0775, Ff0775, Mf0775, Tf0775, Ag0775, Hg0775, Og0775, Vg0775, Ch0775, Jh0775;
wire Qh0775, Xh0775, Ei0775, Li0775, Si0775, Zi0775, Gj0775, Nj0775, Uj0775, Bk0775;
wire Ik0775, Pk0775, Wk0775, Dl0775, Kl0775, Rl0775, Yl0775, Fm0775, Mm0775, Tm0775;
wire An0775, Hn0775, On0775, Vn0775, Co0775, Jo0775, Qo0775, Xo0775, Ep0775, Lp0775;
wire Sp0775, Zp0775, Gq0775, Nq0775, Uq0775, Br0775, Ir0775, Pr0775, Wr0775, Ds0775;
wire Ks0775, Rs0775, Ys0775, Ft0775, Mt0775, Tt0775, Au0775, Hu0775, Ou0775, Vu0775;
wire Cv0775, Jv0775, Qv0775, Xv0775, Ew0775, Lw0775, Sw0775, Zw0775, Gx0775, Nx0775;
wire Ux0775, By0775, Iy0775, Py0775, Wy0775, Dz0775, Kz0775, Rz0775, Yz0775, F01775;
wire M01775, T01775, A11775, H11775, O11775, V11775, C21775, J21775, Q21775, X21775;
wire E31775, L31775, S31775, Z31775, G41775, N41775, U41775, B51775, I51775, P51775;
wire W51775, D61775, K61775, R61775, Y61775, F71775, M71775, T71775, A81775, H81775;
wire O81775, V81775, C91775, J91775, Q91775, X91775, Ea1775, La1775, Sa1775, Za1775;
wire Gb1775, Nb1775, Ub1775, Bc1775, Ic1775, Pc1775, Wc1775, Dd1775, Kd1775, Rd1775;
wire Yd1775, Fe1775, Me1775, Te1775, Af1775, Hf1775, Of1775, Vf1775, Cg1775, Jg1775;
wire Qg1775, Xg1775, Eh1775, Lh1775, Sh1775, Zh1775, Gi1775, Ni1775, Ui1775, Bj1775;
wire Ij1775, Pj1775, Wj1775, Dk1775, Kk1775, Rk1775, Yk1775, Fl1775, Ml1775, Tl1775;
wire Am1775, Hm1775, Om1775, Vm1775, Cn1775, Jn1775, Qn1775, Xn1775, Eo1775, Lo1775;
wire So1775, Zo1775, Gp1775, Np1775, Up1775, Bq1775, Iq1775, Pq1775, Wq1775, Dr1775;
wire Kr1775, Rr1775, Yr1775, Fs1775, Ms1775, Ts1775, At1775, Ht1775, Ot1775, Vt1775;
wire Cu1775, Ju1775, Qu1775, Xu1775, Ev1775, Lv1775, Sv1775, Zv1775, Gw1775, Nw1775;
wire Uw1775, Bx1775, Ix1775, Px1775, Wx1775, Dy1775, Ky1775, Ry1775, Yy1775, Fz1775;
wire Mz1775, Tz1775, A02775, H02775, O02775, V02775, C12775, J12775, Q12775, X12775;
wire E22775, L22775, S22775, Z22775, G32775, N32775, U32775, B42775, I42775, P42775;
wire W42775, D52775, K52775, R52775, Y52775, F62775, M62775, T62775, A72775, H72775;
wire O72775, V72775, C82775, J82775, Q82775, X82775, E92775, L92775, S92775, Z92775;
wire Ga2775, Na2775, Ua2775, Bb2775, Ib2775, Pb2775, Wb2775, Dc2775, Kc2775, Rc2775;
wire Yc2775, Fd2775, Md2775, Td2775, Ae2775, He2775, Oe2775, Ve2775, Cf2775, Jf2775;
wire Qf2775, Xf2775, Eg2775, Lg2775, Sg2775, Zg2775, Gh2775, Nh2775, Uh2775, Bi2775;
wire Ii2775, Pi2775, Wi2775, Dj2775, Kj2775, Rj2775, Yj2775, Fk2775, Mk2775, Tk2775;
wire Al2775, Hl2775, Ol2775, Vl2775, Cm2775, Jm2775, Qm2775, Xm2775, En2775, Ln2775;
wire Sn2775, Zn2775, Go2775, No2775, Uo2775, Bp2775, Ip2775, Pp2775, Wp2775, Dq2775;
wire Kq2775, Rq2775, Yq2775, Fr2775, Mr2775, Tr2775, As2775, Hs2775, Os2775, Vs2775;
wire Ct2775, Jt2775, Qt2775, Xt2775, Eu2775, Lu2775, Su2775, Zu2775, Gv2775, Nv2775;
wire Uv2775, Bw2775, Iw2775, Pw2775, Ww2775, Dx2775, Kx2775, Rx2775, Yx2775, Fy2775;
wire My2775, Ty2775, Az2775, Hz2775, Oz2775, Vz2775, C03775, J03775, Q03775, X03775;
wire E13775, L13775, S13775, Z13775, G23775, N23775, U23775, B33775, I33775, P33775;
wire W33775, D43775, K43775, R43775, Y43775, F53775, M53775, T53775, A63775, H63775;
wire O63775, V63775, C73775, J73775, Q73775, X73775, E83775, L83775, S83775, Z83775;
wire G93775, N93775, U93775, Ba3775, Ia3775, Pa3775, Wa3775, Db3775, Kb3775, Rb3775;
wire Yb3775, Fc3775, Mc3775, Tc3775, Ad3775, Hd3775, Od3775, Vd3775, Ce3775, Je3775;
wire Qe3775, Xe3775, Ef3775, Lf3775, Sf3775, Zf3775, Gg3775, Ng3775, Ug3775, Bh3775;
wire Ih3775, Ph3775, Wh3775, Di3775, Ki3775, Ri3775, Yi3775, Fj3775, Mj3775, Tj3775;
wire Ak3775, Hk3775, Ok3775, Vk3775, Cl3775, Jl3775, Ql3775, Xl3775, Em3775, Lm3775;
wire Sm3775, Zm3775, Gn3775, Nn3775, Un3775, Bo3775, Io3775, Po3775, Wo3775, Dp3775;
wire Kp3775, Rp3775, Yp3775, Fq3775, Mq3775, Tq3775, Ar3775, Hr3775, Or3775, Vr3775;
wire Cs3775, Js3775, Qs3775, Xs3775, Et3775, Lt3775, St3775, Zt3775, Gu3775, Nu3775;
wire Uu3775, Bv3775, Iv3775, Pv3775, Wv3775, Dw3775, Kw3775, Rw3775, Yw3775, Fx3775;
wire Mx3775, Tx3775, Ay3775, Hy3775, Oy3775, Vy3775, Cz3775, Jz3775, Qz3775, Xz3775;
wire E04775, L04775, S04775, Z04775, G14775, N14775, U14775, B24775, I24775, P24775;
wire W24775, D34775, K34775, R34775, Y34775, F44775, M44775, T44775, A54775, H54775;
wire O54775, V54775, C64775, J64775, Q64775, X64775, E74775, L74775, S74775, Z74775;
wire G84775, N84775, U84775, B94775, I94775, P94775, W94775, Da4775, Ka4775, Ra4775;
wire Ya4775, Fb4775, Mb4775, Tb4775, Ac4775, Hc4775, Oc4775, Vc4775, Cd4775, Jd4775;
wire Qd4775, Xd4775, Ee4775, Le4775, Se4775, Ze4775, Gf4775, Nf4775, Uf4775, Bg4775;
wire Ig4775, Pg4775, Wg4775, Dh4775, Kh4775, Rh4775, Yh4775, Fi4775, Mi4775, Ti4775;
wire Aj4775, Hj4775, Oj4775, Vj4775, Ck4775, Jk4775, Qk4775, Xk4775, El4775, Ll4775;
wire Sl4775, Zl4775, Gm4775, Nm4775, Um4775, Bn4775, In4775, Pn4775, Wn4775, Do4775;
wire Ko4775, Ro4775, Yo4775, Fp4775, Mp4775, Tp4775, Aq4775, Hq4775, Oq4775, Vq4775;
wire Cr4775, Jr4775, Qr4775, Xr4775, Es4775, Ls4775, Ss4775, Zs4775, Gt4775, Nt4775;
wire Ut4775, Bu4775, Iu4775, Pu4775, Wu4775, Dv4775, Kv4775, Rv4775, Yv4775, Fw4775;
wire Mw4775, Tw4775, Ax4775, Hx4775, Ox4775, Vx4775, Cy4775, Jy4775, Qy4775, Xy4775;
wire Ez4775, Lz4775, Sz4775, Zz4775, G05775, N05775, U05775, B15775, I15775, P15775;
wire W15775, D25775, K25775, R25775, Y25775, F35775, M35775, T35775, A45775, H45775;
wire O45775, V45775, C55775, J55775, Q55775, X55775, E65775, L65775, S65775, Z65775;
wire G75775, N75775, U75775, B85775, I85775, P85775, W85775, D95775, K95775, R95775;
wire Y95775, Fa5775, Ma5775, Ta5775, Ab5775, Hb5775, Ob5775, Vb5775, Cc5775, Jc5775;
wire Qc5775, Xc5775, Ed5775, Ld5775, Sd5775, Zd5775, Ge5775, Ne5775, Ue5775, Bf5775;
wire If5775, Pf5775, Wf5775, Dg5775, Kg5775, Rg5775, Yg5775, Fh5775, Mh5775, Th5775;
wire Ai5775, Hi5775, Oi5775, Vi5775, Cj5775, Jj5775, Qj5775, Xj5775, Ek5775, Lk5775;
wire Sk5775, Zk5775, Gl5775, Nl5775, Ul5775, Bm5775, Im5775, Pm5775, Wm5775, Dn5775;
wire Kn5775, Rn5775, Yn5775, Fo5775, Mo5775, To5775, Ap5775, Hp5775, Op5775, Vp5775;
wire Cq5775, Jq5775, Qq5775, Xq5775, Er5775, Lr5775, Sr5775, Zr5775, Gs5775, Ns5775;
wire Us5775, Bt5775, It5775, Pt5775, Wt5775, Du5775, Ku5775, Ru5775, Yu5775, Fv5775;
wire Mv5775, Tv5775, Aw5775, Hw5775, Ow5775, Vw5775, Cx5775, Jx5775, Qx5775, Xx5775;
wire Ey5775, Ly5775, Sy5775, Zy5775, Gz5775, Nz5775, Uz5775, B06775, I06775, P06775;
wire W06775, D16775, K16775, R16775, Y16775, F26775, M26775, T26775, A36775, H36775;
wire O36775, V36775, C46775, J46775, Q46775, X46775, E56775, L56775, S56775, Z56775;
wire G66775, N66775, U66775, B76775, I76775, P76775, W76775, D86775, K86775, R86775;
wire Y86775, F96775, M96775, T96775, Aa6775, Ha6775, Oa6775, Va6775, Cb6775, Jb6775;
wire Qb6775, Xb6775, Ec6775, Lc6775, Sc6775, Zc6775, Gd6775, Nd6775, Ud6775, Be6775;
wire Ie6775, Pe6775, We6775, Df6775, Kf6775, Rf6775, Yf6775, Fg6775, Mg6775, Tg6775;
wire Ah6775, Hh6775, Oh6775, Vh6775, Ci6775, Ji6775, Qi6775, Xi6775, Ej6775, Lj6775;
wire Sj6775, Zj6775, Gk6775, Nk6775, Uk6775, Bl6775, Il6775, Pl6775, Wl6775, Dm6775;
wire Km6775, Rm6775, Ym6775, Fn6775, Mn6775, Tn6775, Ao6775, Ho6775, Oo6775, Vo6775;
wire Cp6775, Jp6775, Qp6775, Xp6775, Eq6775, Lq6775, Sq6775, Zq6775, Gr6775, Nr6775;
wire Ur6775, Bs6775, Is6775, Ps6775, Ws6775, Dt6775, Kt6775, Rt6775, Yt6775, Fu6775;
wire Mu6775, Tu6775, Av6775, Hv6775, Ov6775, Vv6775, Cw6775, Jw6775, Qw6775, Xw6775;
wire Ex6775, Lx6775, Sx6775, Zx6775, Gy6775, Ny6775, Uy6775, Bz6775, Iz6775, Pz6775;
wire Wz6775, D07775, K07775, R07775, Y07775, F17775, M17775, T17775, A27775, H27775;
wire O27775, V27775, C37775, J37775, Q37775, X37775, E47775, L47775, S47775, Z47775;
wire G57775, N57775, U57775, B67775, I67775, P67775, W67775, D77775, K77775, R77775;
wire Y77775, F87775, M87775, T87775, A97775, H97775, O97775, V97775, Ca7775, Ja7775;
wire Qa7775, Xa7775, Eb7775, Lb7775, Sb7775, Zb7775, Gc7775, Nc7775, Uc7775, Bd7775;
wire Id7775, Pd7775, Wd7775, De7775, Ke7775, Re7775, Ye7775, Ff7775, Mf7775, Tf7775;
wire Ag7775, Hg7775, Og7775, Vg7775, Ch7775, Jh7775, Qh7775, Xh7775, Ei7775, Li7775;
wire Si7775, Zi7775, Gj7775, Nj7775, Uj7775, Bk7775, Ik7775, Pk7775, Wk7775, Dl7775;
wire Kl7775, Rl7775, Yl7775, Fm7775, Mm7775, Tm7775, An7775, Hn7775, On7775, Vn7775;
wire Co7775, Jo7775, Qo7775, Xo7775, Ep7775, Lp7775, Sp7775, Zp7775, Gq7775, Nq7775;
wire Uq7775, Br7775, Ir7775, Pr7775, Wr7775, Ds7775, Ks7775, Rs7775, Ys7775, Ft7775;
wire Mt7775, Tt7775, Au7775, Hu7775, Ou7775, Vu7775, Cv7775, Jv7775, Qv7775, Xv7775;
wire Ew7775, Lw7775, Sw7775, Zw7775, Gx7775, Nx7775, Ux7775, By7775, Iy7775, Py7775;
wire Wy7775, Dz7775, Kz7775, Rz7775, Yz7775, F08775, M08775, T08775, A18775, H18775;
wire O18775, V18775, C28775, J28775, Q28775, X28775, E38775, L38775, S38775, Z38775;
wire G48775, N48775, U48775, B58775, I58775, P58775, W58775, D68775, K68775, R68775;
wire Y68775, F78775, M78775, T78775, A88775, H88775, O88775, V88775, C98775, J98775;
wire Q98775, X98775, Ea8775, La8775, Sa8775, Za8775, Gb8775, Nb8775, Ub8775, Bc8775;
wire Ic8775, Pc8775, Wc8775, Dd8775, Kd8775, Rd8775, Yd8775, Fe8775, Me8775, Te8775;
wire Af8775, Hf8775, Of8775, Vf8775, Cg8775, Jg8775, Qg8775, Xg8775, Eh8775, Lh8775;
wire Sh8775, Zh8775, Gi8775, Ni8775, Ui8775, Bj8775, Ij8775, Pj8775, Wj8775, Dk8775;
wire Kk8775, Rk8775, Yk8775, Fl8775, Ml8775, Tl8775, Am8775, Hm8775, Om8775, Vm8775;
wire Cn8775, Jn8775, Qn8775, Xn8775, Eo8775, Lo8775, So8775, Zo8775, Gp8775, Np8775;
wire Up8775, Bq8775, Iq8775, Pq8775, Wq8775, Dr8775, Kr8775, Rr8775, Yr8775, Fs8775;
wire Ms8775, Ts8775, At8775, Ht8775, Ot8775, Vt8775, Cu8775, Ju8775, Qu8775, Xu8775;
wire Ev8775, Lv8775, Sv8775, Zv8775, Gw8775, Nw8775, Uw8775, Bx8775, Ix8775, Px8775;
wire Wx8775, Dy8775, Ky8775, Ry8775, Yy8775, Fz8775, Mz8775, Tz8775, A09775, H09775;
wire O09775, V09775, C19775, J19775, Q19775, X19775, E29775, L29775, S29775, Z29775;
wire G39775, N39775, U39775, B49775, I49775, P49775, W49775, D59775, K59775, R59775;
wire Y59775, F69775, M69775, T69775, A79775, H79775, O79775, V79775, C89775, J89775;
wire Q89775, X89775, E99775, L99775, S99775, Z99775, Ga9775, Na9775, Ua9775, Bb9775;
wire Ib9775, Pb9775, Wb9775, Dc9775, Kc9775, Rc9775, Yc9775, Fd9775, Md9775, Td9775;
wire Ae9775, He9775, Oe9775, Ve9775, Cf9775, Jf9775, Qf9775, Xf9775, Eg9775, Lg9775;
wire Sg9775, Zg9775, Gh9775, Nh9775, Uh9775, Bi9775, Ii9775, Pi9775, Wi9775, Dj9775;
wire Kj9775, Rj9775, Yj9775, Fk9775, Mk9775, Tk9775, Al9775, Hl9775, Ol9775, Vl9775;
wire Cm9775, Jm9775, Qm9775, Xm9775, En9775, Ln9775, Sn9775, Zn9775, Go9775, No9775;
wire Uo9775, Bp9775, Ip9775, Pp9775, Wp9775, Dq9775, Kq9775, Rq9775, Yq9775, Fr9775;
wire Mr9775, Tr9775, As9775, Hs9775, Os9775, Vs9775, Ct9775, Jt9775, Qt9775, Xt9775;
wire Eu9775, Lu9775, Su9775, Zu9775, Gv9775, Nv9775, Uv9775, Bw9775, Iw9775, Pw9775;
wire Ww9775, Dx9775, Kx9775, Rx9775, Yx9775, Fy9775, My9775, Ty9775, Az9775, Hz9775;
wire Oz9775, Vz9775, C0a775, J0a775, Q0a775, X0a775, E1a775, L1a775, S1a775, Z1a775;
wire G2a775, N2a775, U2a775, B3a775, I3a775, P3a775, W3a775, D4a775, K4a775, R4a775;
wire Y4a775, F5a775, M5a775, T5a775, A6a775, H6a775, O6a775, V6a775, C7a775, J7a775;
wire Q7a775, X7a775, E8a775, L8a775, S8a775, Z8a775, G9a775, N9a775, U9a775, Baa775;
wire Iaa775, Paa775, Waa775, Dba775, Kba775, Rba775, Yba775, Fca775, Mca775, Tca775;
wire Ada775, Hda775, Oda775, Vda775, Cea775, Jea775, Qea775, Xea775, Efa775, Lfa775;
wire Sfa775, Zfa775, Gga775, Nga775, Uga775, Bha775, Iha775, Pha775, Wha775, Dia775;
wire Kia775, Ria775, Yia775, Fja775, Mja775, Tja775, Aka775, Hka775, Oka775, Vka775;
wire Cla775, Jla775, Qla775, Xla775, Ema775, Lma775, Sma775, Zma775, Gna775, Nna775;
wire Una775, Boa775, Ioa775, Poa775, Woa775, Dpa775, Kpa775, Rpa775, Ypa775, Fqa775;
wire Mqa775, Tqa775, Ara775, Hra775, Ora775, Vra775, Csa775, Jsa775, Qsa775, Xsa775;
wire Eta775, Lta775, Sta775, Zta775, Gua775, Nua775, Uua775, Bva775, Iva775, Pva775;
wire Wva775, Dwa775, Kwa775, Rwa775, Ywa775, Fxa775, Mxa775, Txa775, Aya775, Hya775;
wire Oya775, Vya775, Cza775, Jza775, Qza775, Xza775, E0b775, L0b775, S0b775, Z0b775;
wire G1b775, N1b775, U1b775, B2b775, I2b775, P2b775, W2b775, D3b775, K3b775, R3b775;
wire Y3b775, F4b775, M4b775, T4b775, A5b775, H5b775, O5b775, V5b775, C6b775, J6b775;
wire Q6b775, X6b775, E7b775, L7b775, S7b775, Z7b775, G8b775, N8b775, U8b775, B9b775;
wire I9b775, P9b775, W9b775, Dab775, Kab775, Rab775, Yab775, Fbb775, Mbb775, Tbb775;
wire Acb775, Hcb775, Ocb775, Vcb775, Cdb775, Jdb775, Qdb775, Xdb775, Eeb775, Leb775;
wire Seb775, Zeb775, Gfb775, Nfb775, Ufb775, Bgb775, Igb775, Pgb775, Wgb775, Dhb775;
wire Khb775, Rhb775, Yhb775, Fib775, Mib775, Tib775, Ajb775, Hjb775, Ojb775, Vjb775;
wire Ckb775, Jkb775, Qkb775, Xkb775, Elb775, Llb775, Slb775, Zlb775, Gmb775, Nmb775;
wire Umb775, Bnb775, Inb775, Pnb775, Wnb775, Dob775, Kob775, Rob775, Yob775, Fpb775;
wire Mpb775, Tpb775, Aqb775, Hqb775, Oqb775, Vqb775, Crb775, Jrb775, Qrb775, Xrb775;
wire Esb775, Lsb775, Ssb775, Zsb775, Gtb775, Ntb775, Utb775, Bub775, Iub775, Pub775;
wire Wub775, Dvb775, Kvb775, Rvb775, Yvb775, Fwb775, Mwb775, Twb775, Axb775, Hxb775;
wire Oxb775, Vxb775, Cyb775, Jyb775, Qyb775, Xyb775, Ezb775, Lzb775, Szb775, Zzb775;
wire G0c775, N0c775, U0c775, B1c775, I1c775, P1c775, W1c775, D2c775, K2c775, R2c775;
wire Y2c775, F3c775, M3c775, T3c775, A4c775, H4c775, O4c775, V4c775, C5c775, J5c775;
wire Q5c775, X5c775, E6c775, L6c775, S6c775, Z6c775, G7c775, N7c775, U7c775, B8c775;
wire I8c775, P8c775, W8c775, D9c775, K9c775, R9c775, Y9c775, Fac775, Mac775, Tac775;
wire Abc775, Hbc775, Obc775, Vbc775, Ccc775, Jcc775, Qcc775, Xcc775, Edc775, Ldc775;
wire Sdc775, Zdc775, Gec775, Nec775, Uec775, Bfc775, Ifc775, Pfc775, Wfc775, Dgc775;
wire Kgc775, Rgc775, Ygc775, Fhc775, Mhc775, Thc775, Aic775, Hic775, Oic775, Vic775;
wire Cjc775, Jjc775, Qjc775, Xjc775, Ekc775, Lkc775, Skc775, Zkc775, Glc775, Nlc775;
wire Ulc775, Bmc775, Imc775, Pmc775, Wmc775, Dnc775, Knc775, Rnc775, Ync775, Foc775;
wire Moc775, Toc775, Apc775, Hpc775, Opc775, Vpc775, Cqc775, Jqc775, Qqc775, Xqc775;
wire Erc775, Lrc775, Src775, Zrc775, Gsc775, Nsc775, Usc775, Btc775, Itc775, Ptc775;
wire Wtc775, Duc775, Kuc775, Ruc775, Yuc775, Fvc775, Mvc775, Tvc775, Awc775, Hwc775;
wire Owc775, Vwc775, Cxc775, Jxc775, Qxc775, Xxc775, Eyc775, Lyc775, Syc775, Zyc775;
wire Gzc775, Nzc775, Uzc775, B0d775, I0d775, P0d775, W0d775, D1d775, K1d775, R1d775;
wire Y1d775, F2d775, M2d775, T2d775, A3d775, H3d775, O3d775, V3d775, C4d775, J4d775;
wire Q4d775, X4d775, E5d775, L5d775, S5d775, Z5d775, G6d775, N6d775, U6d775, B7d775;
wire I7d775, P7d775, W7d775, D8d775, K8d775, R8d775, Y8d775, F9d775, M9d775, T9d775;
wire Aad775, Had775, Oad775, Vad775, Cbd775, Jbd775, Qbd775, Xbd775, Ecd775, Lcd775;
wire Scd775, Zcd775, Gdd775, Ndd775, Udd775, Bed775, Ied775, Ped775, Wed775, Dfd775;
wire Kfd775, Rfd775, Yfd775, Fgd775, Mgd775, Tgd775, Ahd775, Hhd775, Ohd775, Vhd775;
wire Cid775, Jid775, Qid775, Xid775, Ejd775, Ljd775, Sjd775, Zjd775, Gkd775, Nkd775;
wire Ukd775, Bld775, Ild775, Pld775, Wld775, Dmd775, Kmd775, Rmd775, Ymd775, Fnd775;
wire Mnd775, Tnd775, Aod775, Hod775, Ood775, Vod775, Cpd775, Jpd775, Qpd775, Xpd775;
wire Eqd775, Lqd775, Sqd775, Zqd775, Grd775, Nrd775, Urd775, Bsd775, Isd775, Psd775;
wire Wsd775, Dtd775, Ktd775, Rtd775, Ytd775, Fud775, Mud775, Tud775, Avd775, Hvd775;
wire Ovd775, Vvd775, Cwd775, Jwd775, Qwd775, Xwd775, Exd775, Lxd775, Sxd775, Zxd775;
wire Gyd775, Nyd775, Uyd775, Bzd775, Izd775, Pzd775, Wzd775, D0e775, K0e775, R0e775;
wire Y0e775, F1e775, M1e775, T1e775, A2e775, H2e775, O2e775, V2e775, C3e775, J3e775;
wire Q3e775, X3e775, E4e775, L4e775, S4e775, Z4e775, G5e775, N5e775, U5e775, B6e775;
wire I6e775, P6e775, W6e775, D7e775, K7e775, R7e775, Y7e775, F8e775, M8e775, T8e775;
wire A9e775, H9e775, O9e775, V9e775, Cae775, Jae775, Qae775, Xae775, Ebe775, Lbe775;
wire Sbe775, Zbe775, Gce775, Nce775, Uce775, Bde775, Ide775, Pde775, Wde775, Dee775;
wire Kee775, Ree775, Yee775, Ffe775, Mfe775, Tfe775, Age775, Hge775, Oge775, Vge775;
wire Che775, Jhe775, Qhe775, Xhe775, Eie775, Lie775, Sie775, Zie775, Gje775, Nje775;
wire Uje775, Bke775, Ike775, Pke775, Wke775, Dle775, Kle775, Rle775, Yle775, Fme775;
wire Mme775, Tme775, Ane775, Hne775, One775, Vne775, Coe775, Joe775, Qoe775, Xoe775;
wire Epe775, Lpe775, Spe775, Zpe775, Gqe775, Nqe775, Uqe775, Bre775, Ire775, Pre775;
wire Wre775, Dse775, Kse775, Rse775, Yse775, Fte775, Mte775, Tte775, Aue775, Hue775;
wire Oue775, Vue775, Cve775, Jve775, Qve775, Xve775, Ewe775, Lwe775, Swe775, Zwe775;
wire Gxe775, Nxe775, Uxe775, Bye775, Iye775, Pye775, Wye775, Dze775, Kze775, Rze775;
wire Yze775, F0f775, M0f775, T0f775, A1f775, H1f775, O1f775, V1f775, C2f775, J2f775;
wire Q2f775, X2f775, E3f775, L3f775, S3f775, Z3f775, G4f775, N4f775, U4f775, B5f775;
wire I5f775, P5f775, W5f775, D6f775, K6f775, R6f775, Y6f775, F7f775, M7f775, T7f775;
wire A8f775, H8f775, O8f775, V8f775, C9f775, J9f775, Q9f775, X9f775, Eaf775, Laf775;
wire Saf775, Zaf775, Gbf775, Nbf775, Ubf775, Bcf775, Icf775, Pcf775, Wcf775, Ddf775;
wire Kdf775, Rdf775, Ydf775, Fef775, Mef775, Tef775, Aff775, Hff775, Off775, Vff775;
wire Cgf775, Jgf775, Qgf775, Xgf775, Ehf775, Lhf775, Shf775, Zhf775, Gif775, Nif775;
wire Uif775, Bjf775, Ijf775, Pjf775, Wjf775, Dkf775, Kkf775, Rkf775, Ykf775, Flf775;
wire Mlf775, Tlf775, Amf775, Hmf775, Omf775, Vmf775, Cnf775, Jnf775, Qnf775, Xnf775;
wire Eof775, Lof775, Sof775, Zof775, Gpf775, Npf775, Upf775, Bqf775, Iqf775, Pqf775;
wire Wqf775, Drf775, Krf775, Rrf775, Yrf775, Fsf775, Msf775, Tsf775, Atf775, Htf775;
wire Otf775, Vtf775, Cuf775, Juf775, Quf775, Xuf775, Evf775, Lvf775, Svf775, Zvf775;
wire Gwf775, Nwf775, Uwf775, Bxf775, Ixf775, Pxf775, Wxf775, Dyf775, Kyf775, Ryf775;
wire Yyf775, Fzf775, Mzf775, Tzf775, A0g775, H0g775, O0g775, V0g775, C1g775, J1g775;
wire Q1g775, X1g775, E2g775, L2g775, S2g775, Z2g775, G3g775, N3g775, U3g775, B4g775;
wire I4g775, P4g775, W4g775, D5g775, K5g775, R5g775, Y5g775, F6g775, M6g775, T6g775;
wire A7g775, H7g775, O7g775, V7g775, C8g775, J8g775, Q8g775, X8g775, E9g775, L9g775;
wire S9g775, Z9g775, Gag775, Nag775, Uag775, Bbg775, Ibg775, Pbg775, Wbg775, Dcg775;
wire Kcg775, Rcg775, Ycg775, Fdg775, Mdg775, Tdg775, Aeg775, Heg775, Oeg775, Veg775;
wire Cfg775, Jfg775, Qfg775, Xfg775, Egg775, Lgg775, Sgg775, Zgg775, Ghg775, Nhg775;
wire Uhg775, Big775, Iig775, Pig775, Wig775, Djg775, Kjg775, Rjg775, Yjg775, Fkg775;
wire Mkg775, Tkg775, Alg775, Hlg775, Olg775, Vlg775, Cmg775, Jmg775, Qmg775, Xmg775;
wire Eng775, Lng775, Sng775, Zng775, Gog775, Nog775, Uog775, Bpg775, Ipg775, Ppg775;
wire Wpg775, Dqg775, Kqg775, Rqg775, Yqg775, Frg775, Mrg775, Trg775, Asg775, Hsg775;
wire Osg775, Vsg775, Ctg775, Jtg775, Qtg775, Xtg775, Eug775, Lug775, Sug775, Zug775;
wire Gvg775, Nvg775, Uvg775, Bwg775, Iwg775, Pwg775, Wwg775, Dxg775, Kxg775, Rxg775;
wire Yxg775, Fyg775, Myg775, Tyg775, Azg775, Hzg775, Ozg775, Vzg775, C0h775, J0h775;
wire Q0h775, X0h775, E1h775, L1h775, S1h775, Z1h775, G2h775, N2h775, U2h775, B3h775;
wire I3h775, P3h775, W3h775, D4h775, K4h775, R4h775, Y4h775, F5h775, M5h775, T5h775;
wire A6h775, H6h775, O6h775, V6h775, C7h775, J7h775, Q7h775, X7h775, E8h775, L8h775;
wire S8h775, Z8h775, G9h775, N9h775, U9h775, Bah775, Iah775, Pah775, Wah775, Dbh775;
wire Kbh775, Rbh775, Ybh775, Fch775, Mch775, Tch775, Adh775, Hdh775, Odh775, Vdh775;
wire Ceh775, Jeh775, Qeh775, Xeh775, Efh775, Lfh775, Sfh775, Zfh775, Ggh775, Ngh775;
wire Ugh775, Bhh775, Ihh775, Phh775, Whh775, Dih775, Kih775, Rih775, Yih775, Fjh775;
wire Mjh775, Tjh775, Akh775, Hkh775, Okh775, Vkh775, Clh775, Jlh775, Qlh775, Xlh775;
wire Emh775, Lmh775, Smh775, Zmh775, Gnh775, Nnh775, Unh775, Boh775, Ioh775, Poh775;
wire Woh775, Dph775, Kph775, Rph775, Yph775, Fqh775, Mqh775, Tqh775, Arh775, Hrh775;
wire Orh775, Vrh775, Csh775, Jsh775, Qsh775, Xsh775, Eth775, Lth775, Sth775, Zth775;
wire Guh775, Nuh775, Uuh775, Bvh775, Ivh775, Pvh775, Wvh775, Dwh775, Kwh775, Rwh775;
wire Ywh775, Fxh775, Mxh775, Txh775, Ayh775, Hyh775, Oyh775, Vyh775, Czh775, Jzh775;
wire Qzh775, Xzh775, E0i775, L0i775, S0i775, Z0i775, G1i775, N1i775, U1i775, B2i775;
wire I2i775, P2i775, W2i775, D3i775, K3i775, R3i775, Y3i775, F4i775, M4i775, T4i775;
wire A5i775, H5i775, O5i775, V5i775, C6i775, J6i775, Q6i775, X6i775, E7i775, L7i775;
wire S7i775, Z7i775, G8i775, N8i775, U8i775, B9i775, I9i775, P9i775, W9i775, Dai775;
wire Kai775, Rai775, Yai775, Fbi775, Mbi775, Tbi775, Aci775, Hci775, Oci775, Vci775;
wire Cdi775, Jdi775, Qdi775, Xdi775, Eei775, Lei775, Sei775, Zei775, Gfi775, Nfi775;
wire Ufi775, Bgi775, Igi775, Pgi775, Wgi775, Dhi775, Khi775, Rhi775, Yhi775, Fii775;
wire Mii775, Tii775, Aji775, Hji775, Oji775, Vji775, Cki775, Jki775, Qki775, Xki775;
wire Eli775, Lli775, Sli775, Zli775, Gmi775, Nmi775, Umi775, Bni775, Ini775, Pni775;
wire Wni775, Doi775, Koi775, Roi775, Yoi775, Fpi775, Mpi775, Tpi775, Aqi775, Hqi775;
wire Oqi775, Vqi775, Cri775, Jri775, Qri775, Xri775, Esi775, Lsi775, Ssi775, Zsi775;
wire Gti775, Nti775, Uti775, Bui775, Iui775, Pui775, Wui775, Dvi775, Kvi775, Rvi775;
wire Yvi775, Fwi775, Mwi775, Twi775, Axi775, Hxi775, Oxi775, Vxi775, Cyi775, Jyi775;
wire Qyi775, Xyi775, Ezi775, Lzi775, Szi775, Zzi775, G0j775, N0j775, U0j775, B1j775;
wire I1j775, P1j775, W1j775, D2j775, K2j775, R2j775, Y2j775, F3j775, M3j775, T3j775;
wire A4j775, H4j775, O4j775, V4j775, C5j775, J5j775, Q5j775, X5j775, E6j775, L6j775;
wire S6j775, Z6j775, G7j775, N7j775, U7j775, B8j775, I8j775, P8j775, W8j775, D9j775;
wire K9j775, R9j775, Y9j775, Faj775, Maj775, Taj775, Abj775, Hbj775, Obj775, Vbj775;
wire Ccj775, Jcj775, Qcj775, Xcj775, Edj775, Ldj775, Sdj775, Zdj775, Gej775, Nej775;
wire Uej775, Bfj775, Ifj775, Pfj775, Wfj775, Dgj775, Kgj775, Rgj775, Ygj775, Fhj775;
wire Mhj775, Thj775, Aij775, Hij775, Oij775, Vij775, Cjj775, Jjj775, Qjj775, Xjj775;
wire Ekj775, Lkj775, Skj775, Zkj775, Glj775, Nlj775, Ulj775, Bmj775, Imj775, Pmj775;
wire Wmj775, Dnj775, Knj775, Rnj775, Ynj775, Foj775, Moj775, Toj775, Apj775, Hpj775;
wire Opj775, Vpj775, Cqj775, Jqj775, Qqj775, Xqj775, Erj775, Lrj775, Srj775, Zrj775;
wire Gsj775, Nsj775, Usj775, Btj775, Itj775, Ptj775, Wtj775, Duj775, Kuj775, Ruj775;
wire Yuj775, Fvj775, Mvj775, Tvj775, Awj775, Hwj775, Owj775, Vwj775, Cxj775, Jxj775;
wire Qxj775, Xxj775, Eyj775, Lyj775, Syj775, Zyj775, Gzj775, Nzj775, Uzj775, B0k775;
wire I0k775, P0k775, W0k775, D1k775, K1k775, R1k775, Y1k775, F2k775, M2k775, T2k775;
wire A3k775, H3k775, O3k775, V3k775, C4k775, J4k775, Q4k775, X4k775, E5k775, L5k775;
wire S5k775, Z5k775, G6k775, N6k775, U6k775, B7k775, I7k775, P7k775, W7k775, D8k775;
wire K8k775, R8k775, Y8k775, F9k775, M9k775, T9k775, Aak775, Hak775, Oak775, Vak775;
wire Cbk775, Jbk775, Qbk775, Xbk775, Eck775, Lck775, Sck775, Zck775, Gdk775, Ndk775;
wire Udk775, Bek775, Iek775, Pek775, Wek775, Dfk775, Kfk775, Rfk775, Yfk775, Fgk775;
wire Mgk775, Tgk775, Ahk775, Hhk775, Ohk775, Vhk775, Cik775, Jik775, Qik775, Xik775;
wire Ejk775, Ljk775, Sjk775, Zjk775, Gkk775, Nkk775, Ukk775, Blk775, Ilk775, Plk775;
wire Wlk775, Dmk775, Kmk775, Rmk775, Ymk775, Fnk775, Mnk775, Tnk775, Aok775, Hok775;
wire Ook775, Vok775, Cpk775, Jpk775, Qpk775, Xpk775, Eqk775, Lqk775, Sqk775, Zqk775;
wire Grk775, Nrk775, Urk775, Bsk775, Isk775, Psk775, Wsk775, Dtk775, Ktk775, Rtk775;
wire Ytk775, Fuk775, Muk775, Tuk775, Avk775, Hvk775, Ovk775, Vvk775, Cwk775, Jwk775;
wire Qwk775, Xwk775, Exk775, Lxk775, Sxk775, Zxk775, Gyk775, Nyk775, Uyk775, Bzk775;
wire Izk775, Pzk775, Wzk775, D0l775, K0l775, R0l775, Y0l775, F1l775, M1l775, T1l775;
wire A2l775, H2l775, O2l775, V2l775, C3l775, J3l775, Q3l775, X3l775, E4l775, L4l775;
wire S4l775, Z4l775, G5l775, N5l775, U5l775, B6l775, I6l775, P6l775, W6l775, D7l775;
wire K7l775, R7l775, Y7l775, F8l775, M8l775, T8l775, A9l775, H9l775, O9l775, V9l775;
wire Cal775, Jal775, Qal775, Xal775, Ebl775, Lbl775, Sbl775, Zbl775, Gcl775, Ncl775;
wire Ucl775, Bdl775, Idl775, Pdl775, Wdl775, Del775, Kel775, Rel775, Yel775, Ffl775;
wire Mfl775, Tfl775, Agl775, Hgl775, Ogl775, Vgl775, Chl775, Jhl775, Qhl775, Xhl775;
wire Eil775, Lil775, Sil775, Zil775, Gjl775, Njl775, Ujl775, Bkl775, Ikl775, Pkl775;
wire Wkl775, Dll775, Kll775, Rll775, Yll775, Fml775, Mml775, Tml775, Anl775, Hnl775;
wire Onl775, Vnl775, Col775, Jol775, Qol775, Xol775, Epl775, Lpl775, Spl775, Zpl775;
wire Gql775, Nql775, Uql775, Brl775, Irl775, Prl775, Wrl775, Dsl775, Ksl775, Rsl775;
wire Ysl775, Ftl775, Mtl775, Ttl775, Aul775, Hul775, Oul775, Vul775, Cvl775, Jvl775;
wire Qvl775, Xvl775, Ewl775, Lwl775, Swl775, Zwl775, Gxl775, Nxl775, Uxl775, Byl775;
wire Iyl775, Pyl775, Wyl775, Dzl775, Kzl775, Rzl775, Yzl775, F0m775, M0m775, T0m775;
wire A1m775, H1m775, O1m775, V1m775, C2m775, J2m775, Q2m775, X2m775, E3m775, L3m775;
wire S3m775, Z3m775, G4m775, N4m775, U4m775, B5m775, I5m775, P5m775, W5m775, D6m775;
wire K6m775, R6m775, Y6m775, F7m775, M7m775, T7m775, A8m775, H8m775, O8m775, V8m775;
wire C9m775, J9m775, Q9m775, X9m775, Eam775, Lam775, Sam775, Zam775, Gbm775, Nbm775;
wire Ubm775, Bcm775, Icm775, Pcm775, Wcm775, Ddm775, Kdm775, Rdm775, Ydm775, Fem775;
wire Mem775, Tem775, Afm775, Hfm775, Ofm775, Vfm775, Cgm775, Jgm775, Qgm775, Xgm775;
wire Ehm775, Lhm775, Shm775, Zhm775, Gim775, Nim775, Uim775, Bjm775, Ijm775, Pjm775;
wire Wjm775, Dkm775, Kkm775, Rkm775, Ykm775, Flm775, Mlm775, Tlm775, Amm775, Hmm775;
wire Omm775, Vmm775, Cnm775, Jnm775, Qnm775, Xnm775, Eom775, Lom775, Som775, Zom775;
wire Gpm775, Npm775, Upm775, Bqm775, Iqm775, Pqm775, Wqm775, Drm775, Krm775, Rrm775;
wire Yrm775, Fsm775, Msm775, Tsm775, Atm775, Htm775, Otm775, Vtm775, Cum775, Jum775;
wire Qum775, Xum775, Evm775, Lvm775, Svm775, Zvm775, Gwm775, Nwm775, Uwm775, Bxm775;
wire Ixm775, Pxm775, Wxm775, Dym775, Kym775, Rym775, Yym775, Fzm775, Mzm775, Tzm775;
wire A0n775, H0n775, O0n775, V0n775, C1n775, J1n775, Q1n775, X1n775, E2n775, L2n775;
wire S2n775, Z2n775, G3n775, N3n775, U3n775, B4n775, I4n775, P4n775, W4n775, D5n775;
wire K5n775, R5n775, Y5n775, F6n775, M6n775, T6n775, A7n775, H7n775, O7n775, V7n775;
wire C8n775, J8n775, Q8n775, X8n775, E9n775, L9n775, S9n775, Z9n775, Gan775, Nan775;
wire Uan775, Bbn775, Ibn775, Pbn775, Wbn775, Dcn775, Kcn775, Rcn775, Ycn775, Fdn775;
wire Mdn775, Tdn775, Aen775, Hen775, Oen775, Ven775, Cfn775, Jfn775, Qfn775, Xfn775;
wire Egn775, Lgn775, Sgn775, Zgn775, Ghn775, Nhn775, Uhn775, Bin775, Iin775, Pin775;
wire Win775, Djn775, Kjn775, Rjn775, Yjn775, Fkn775, Mkn775, Tkn775, Aln775, Hln775;
wire Oln775, Vln775, Cmn775, Jmn775, Qmn775, Xmn775, Enn775, Lnn775, Snn775, Znn775;
wire Gon775, Non775, Uon775, Bpn775, Ipn775, Ppn775, Wpn775, Dqn775, Kqn775, Rqn775;
wire Yqn775, Frn775, Mrn775, Trn775, Asn775, Hsn775, Osn775, Vsn775, Ctn775, Jtn775;
wire Qtn775, Xtn775, Eun775, Lun775, Sun775, Zun775, Gvn775, Nvn775, Uvn775, Bwn775;
wire Iwn775, Pwn775, Wwn775, Dxn775, Kxn775, Rxn775, Yxn775, Fyn775, Myn775, Tyn775;
wire Azn775, Hzn775, Ozn775, Vzn775, C0o775, J0o775, Q0o775, X0o775, E1o775, L1o775;
wire S1o775, Z1o775, G2o775, N2o775, U2o775, B3o775, I3o775, P3o775, W3o775, D4o775;
wire K4o775, R4o775, Y4o775, F5o775, M5o775, T5o775, A6o775, H6o775, O6o775, V6o775;
wire C7o775, J7o775, Q7o775, X7o775, E8o775, L8o775, S8o775, Z8o775, G9o775, N9o775;
wire U9o775, Bao775, Iao775, Pao775, Wao775, Dbo775, Kbo775, Rbo775, Ybo775, Fco775;
wire Mco775, Tco775, Ado775, Hdo775, Odo775, Vdo775, Ceo775, Jeo775, Qeo775, Xeo775;
wire Efo775, Lfo775, Sfo775, Zfo775, Ggo775, Ngo775, Ugo775, Bho775, Iho775, Pho775;
wire Who775, Dio775, Kio775, Rio775, Yio775, Fjo775, Mjo775, Tjo775, Ako775, Hko775;
wire Oko775, Vko775, Clo775, Jlo775, Qlo775, Xlo775, Emo775, Lmo775, Smo775, Zmo775;
wire Gno775, Nno775, Uno775, Boo775, Ioo775, Poo775, Woo775, Dpo775, Kpo775, Rpo775;
wire Ypo775, Fqo775, Mqo775, Tqo775, Aro775, Hro775, Oro775, Vro775, Cso775, Jso775;
wire Qso775, Xso775, Eto775, Lto775, Sto775, Zto775, Guo775, Nuo775, Uuo775, Bvo775;
wire Ivo775, Pvo775, Wvo775, Dwo775, Kwo775, Rwo775, Ywo775, Fxo775, Mxo775, Txo775;
wire Ayo775, Hyo775, Oyo775, Vyo775, Czo775, Jzo775, Qzo775, Xzo775, E0p775, L0p775;
wire S0p775, Z0p775, G1p775, N1p775, U1p775, B2p775, I2p775, P2p775, W2p775, D3p775;
wire K3p775, R3p775, Y3p775, F4p775, M4p775, T4p775, A5p775, H5p775, O5p775, V5p775;
wire C6p775, J6p775, Q6p775, X6p775, E7p775, L7p775, S7p775, Z7p775, G8p775, N8p775;
wire U8p775, B9p775, I9p775, P9p775, W9p775, Dap775, Kap775, Rap775, Yap775, Fbp775;
wire Mbp775, Tbp775, Acp775, Hcp775, Ocp775, Vcp775, Cdp775, Jdp775, Qdp775, Xdp775;
wire Eep775, Lep775, Sep775, Zep775, Gfp775, Nfp775, Ufp775, Bgp775, Igp775, Pgp775;
wire Wgp775, Dhp775, Khp775, Rhp775, Yhp775, Fip775, Mip775, Tip775, Ajp775, Hjp775;
wire Ojp775, Vjp775, Ckp775, Jkp775, Qkp775, Xkp775, Elp775, Llp775, Slp775, Zlp775;
wire Gmp775, Nmp775, Ump775, Bnp775, Inp775, Pnp775, Wnp775, Dop775, Kop775, Rop775;
wire Yop775, Fpp775, Mpp775, Tpp775, Aqp775, Hqp775, Oqp775, Vqp775, Crp775, Jrp775;
wire Qrp775, Xrp775, Esp775, Lsp775, Ssp775, Zsp775, Gtp775, Ntp775, Utp775, Bup775;
wire Iup775, Pup775, Wup775, Dvp775, Kvp775, Rvp775, Yvp775, Fwp775, Mwp775, Twp775;
wire Axp775, Hxp775, Oxp775, Vxp775, Cyp775, Jyp775, Qyp775, Xyp775, Ezp775, Lzp775;
wire Szp775, Zzp775, G0q775, N0q775, U0q775, B1q775, I1q775, P1q775, W1q775, D2q775;
wire K2q775, R2q775, Y2q775, F3q775, M3q775, T3q775, A4q775, H4q775, O4q775, V4q775;
wire C5q775, J5q775, Q5q775, X5q775, E6q775, L6q775, S6q775, Z6q775, G7q775, N7q775;
wire U7q775, B8q775, I8q775, P8q775, W8q775, D9q775, K9q775, R9q775, Y9q775, Faq775;
wire Maq775, Taq775, Abq775, Hbq775, Obq775, Vbq775, Ccq775, Jcq775, Qcq775, Xcq775;
wire Edq775, Ldq775, Sdq775, Zdq775, Geq775, Neq775, Ueq775, Bfq775, Ifq775, Pfq775;
wire Wfq775, Dgq775, Kgq775, Rgq775, Ygq775, Fhq775, Mhq775, Thq775, Aiq775, Hiq775;
wire Oiq775, Viq775, Cjq775, Jjq775, Qjq775, Xjq775, Ekq775, Lkq775, Skq775, Zkq775;
wire Glq775, Nlq775, Ulq775, Bmq775, Imq775, Pmq775, Wmq775, Dnq775, Knq775, Rnq775;
wire Ynq775, Foq775, Moq775, Toq775, Apq775, Hpq775, Opq775, Vpq775, Cqq775, Jqq775;
wire Qqq775, Xqq775, Erq775, Lrq775, Srq775, Zrq775, Gsq775, Nsq775, Usq775, Btq775;
wire Itq775, Ptq775, Wtq775, Duq775, Kuq775, Ruq775, Yuq775, Fvq775, Mvq775, Tvq775;
wire Awq775, Hwq775, Owq775, Vwq775, Cxq775, Jxq775, Qxq775, Xxq775, Eyq775, Lyq775;
wire Syq775, Zyq775, Gzq775, Nzq775, Uzq775, B0r775, I0r775, P0r775, W0r775, D1r775;
wire K1r775, R1r775, Y1r775, F2r775, M2r775, T2r775, A3r775, H3r775, O3r775, V3r775;
wire C4r775, J4r775, Q4r775, X4r775, E5r775, L5r775, S5r775, Z5r775, G6r775, N6r775;
wire U6r775, B7r775, I7r775, P7r775, W7r775, D8r775, K8r775, R8r775, Y8r775, F9r775;
wire M9r775, T9r775, Aar775, Har775, Oar775, Var775, Cbr775, Jbr775, Qbr775, Xbr775;
wire Ecr775, Lcr775, Scr775, Zcr775, Gdr775, Ndr775, Udr775, Ber775, Ier775, Per775;
wire Wer775, Dfr775, Kfr775, Rfr775, Yfr775, Fgr775, Mgr775, Tgr775, Ahr775, Hhr775;
wire Ohr775, Vhr775, Cir775, Jir775, Qir775, Xir775, Ejr775, Ljr775, Sjr775, Zjr775;
wire Gkr775, Nkr775, Ukr775, Blr775, Ilr775, Plr775, Wlr775, Dmr775, Kmr775, Rmr775;
wire Ymr775, Fnr775, Mnr775, Tnr775, Aor775, Hor775, Oor775, Vor775, Cpr775, Jpr775;
wire Qpr775, Xpr775, Eqr775, Lqr775, Sqr775, Zqr775, Grr775, Nrr775, Urr775, Bsr775;
wire Isr775, Psr775, Wsr775, Dtr775, Ktr775, Rtr775, Ytr775, Fur775, Mur775, Tur775;
wire Avr775, Hvr775, Ovr775, Vvr775, Cwr775, Jwr775, Qwr775, Xwr775, Exr775, Lxr775;
wire Sxr775, Zxr775, Gyr775, Nyr775, Uyr775, Bzr775, Izr775, Pzr775, Wzr775, D0s775;
wire K0s775, R0s775, Y0s775, F1s775, M1s775, T1s775, A2s775, H2s775, O2s775, V2s775;
wire C3s775, J3s775, Q3s775, X3s775, E4s775, L4s775, S4s775, Z4s775, G5s775, N5s775;
wire U5s775, B6s775, I6s775, P6s775, W6s775, D7s775, K7s775, R7s775, Y7s775, F8s775;
wire M8s775, T8s775, A9s775, H9s775, O9s775, V9s775, Cas775, Jas775, Qas775, Xas775;
wire Ebs775, Lbs775, Sbs775, Zbs775, Gcs775, Ncs775, Ucs775, Bds775, Ids775, Pds775;
wire Wds775, Des775, Kes775, Res775, Yes775, Ffs775, Mfs775, Tfs775, Ags775, Hgs775;
wire Ogs775, Vgs775, Chs775, Jhs775, Qhs775, Xhs775, Eis775, Lis775, Sis775, Zis775;
wire Gjs775, Njs775, Ujs775, Bks775, Iks775, Pks775, Wks775, Dls775, Kls775, Rls775;
wire Yls775, Fms775, Mms775, Tms775, Ans775, Hns775, Ons775, Vns775, Cos775, Jos775;
wire Qos775, Xos775, Eps775, Lps775, Sps775, Zps775, Gqs775, Nqs775, Uqs775, Brs775;
wire Irs775, Prs775, Wrs775, Dss775, Kss775, Rss775, Yss775, Fts775, Mts775, Tts775;
wire Aus775, Hus775, Ous775, Vus775, Cvs775, Jvs775, Qvs775, Xvs775, Ews775, Lws775;
wire Sws775, Zws775, Gxs775, Nxs775, Uxs775, Bys775, Iys775, Pys775, Wys775, Dzs775;
wire Kzs775, Rzs775, Yzs775, F0t775, M0t775, T0t775, A1t775, H1t775, O1t775, V1t775;
wire C2t775, J2t775, Q2t775, X2t775, E3t775, L3t775, S3t775, Z3t775, G4t775, N4t775;
wire U4t775, B5t775, I5t775, P5t775, W5t775, D6t775, K6t775, R6t775, Y6t775, F7t775;
wire M7t775, T7t775, A8t775, H8t775, O8t775, V8t775, C9t775, J9t775, Q9t775, X9t775;
wire Eat775, Lat775, Sat775, Zat775, Gbt775, Nbt775, Ubt775, Bct775, Ict775, Pct775;
wire Wct775, Ddt775, Kdt775, Rdt775, Ydt775, Fet775, Met775, Tet775, Aft775, Hft775;
wire Oft775, Vft775, Cgt775, Jgt775, Qgt775, Xgt775, Eht775, Lht775, Sht775, Zht775;
wire Git775, Nit775, Uit775, Bjt775, Ijt775, Pjt775, Wjt775, Dkt775, Kkt775, Rkt775;
wire Ykt775, Flt775, Mlt775, Tlt775, Amt775, Hmt775, Omt775, Vmt775, Cnt775, Jnt775;
wire Qnt775, Xnt775, Eot775, Lot775, Sot775, Zot775, Gpt775, Npt775, Upt775, Bqt775;
wire Iqt775, Pqt775, Wqt775, Drt775, Krt775, Rrt775, Yrt775, Fst775, Mst775, Tst775;
wire Att775, Htt775, Ott775, Vtt775, Cut775, Jut775, Qut775, Xut775, Evt775, Lvt775;
wire Svt775, Zvt775, Gwt775, Nwt775, Uwt775, Bxt775, Ixt775, Pxt775, Wxt775, Dyt775;
wire Kyt775, Ryt775, Yyt775, Fzt775, Mzt775, Tzt775, A0u775, H0u775, O0u775, V0u775;
wire C1u775, J1u775, Q1u775, X1u775, E2u775, L2u775, S2u775, Z2u775, G3u775, N3u775;
wire U3u775, B4u775, I4u775, P4u775, W4u775, D5u775, K5u775, R5u775, Y5u775, F6u775;
wire M6u775, T6u775, A7u775, H7u775, O7u775, V7u775, C8u775, J8u775, Q8u775, X8u775;
wire E9u775, L9u775, S9u775, Z9u775, Gau775, Nau775, Uau775, Bbu775, Ibu775, Pbu775;
wire Wbu775, Dcu775, Kcu775, Rcu775, Ycu775, Fdu775, Mdu775, Tdu775, Aeu775, Heu775;
wire Oeu775, Veu775, Cfu775, Jfu775, Qfu775, Xfu775, Egu775, Lgu775, Sgu775, Zgu775;
wire Ghu775, Nhu775, Uhu775, Biu775, Iiu775, Piu775, Wiu775, Dju775, Kju775, Rju775;
wire Yju775, Fku775, Mku775, Tku775, Alu775, Hlu775, Olu775, Vlu775, Cmu775, Jmu775;
wire Qmu775, Xmu775, Enu775, Lnu775, Snu775, Znu775, Gou775, Nou775, Uou775, Bpu775;
wire Ipu775, Ppu775, Wpu775, Dqu775, Kqu775, Rqu775, Yqu775, Fru775, Mru775, Tru775;
wire Asu775, Hsu775, Osu775, Vsu775, Ctu775, Jtu775, Qtu775, Xtu775, Euu775, Luu775;
wire Suu775, Zuu775, Gvu775, Nvu775, Uvu775, Bwu775, Iwu775, Pwu775, Wwu775, Dxu775;
wire Kxu775, Rxu775, Yxu775, Fyu775, Myu775, Tyu775, Azu775, Hzu775, Ozu775, Vzu775;
wire C0v775, J0v775, Q0v775, X0v775, E1v775, L1v775, S1v775, Z1v775, G2v775, N2v775;
wire U2v775, B3v775, I3v775, P3v775, W3v775, D4v775, K4v775, R4v775, Y4v775, F5v775;
wire M5v775, T5v775, A6v775, H6v775, O6v775, V6v775, C7v775, J7v775, Q7v775, X7v775;
wire E8v775, L8v775, S8v775, Z8v775, G9v775, N9v775, U9v775, Bav775, Iav775, Pav775;
wire Wav775, Dbv775, Kbv775, Rbv775, Ybv775, Fcv775, Mcv775, Tcv775, Adv775, Hdv775;
wire Odv775, Vdv775, Cev775, Jev775, Qev775, Xev775, Efv775, Lfv775, Sfv775, Zfv775;
wire Ggv775, Ngv775, Ugv775, Bhv775, Ihv775, Phv775, Whv775, Div775, Kiv775, Riv775;
wire Yiv775, Fjv775, Mjv775, Tjv775, Akv775, Hkv775, Okv775, Vkv775, Clv775, Jlv775;
wire Qlv775, Xlv775, Emv775, Lmv775, Smv775, Zmv775, Gnv775, Nnv775, Unv775, Bov775;
wire Iov775, Pov775, Wov775, Dpv775, Kpv775, Rpv775, Ypv775, Fqv775, Mqv775, Tqv775;
wire Arv775, Hrv775, Orv775, Vrv775, Csv775, Jsv775, Qsv775, Xsv775, Etv775, Ltv775;
wire Stv775, Ztv775, Guv775, Nuv775, Uuv775, Bvv775, Ivv775, Pvv775, Wvv775, Dwv775;
wire Kwv775, Rwv775, Ywv775, Fxv775, Mxv775, Txv775, Ayv775, Hyv775, Oyv775, Vyv775;
wire Czv775, Jzv775, Qzv775, Xzv775, E0w775, L0w775, S0w775, Z0w775, G1w775, N1w775;
wire U1w775, B2w775, I2w775, P2w775, W2w775, D3w775, K3w775, R3w775, Y3w775, F4w775;
wire M4w775, T4w775, A5w775, H5w775, O5w775, V5w775, C6w775, J6w775, Q6w775, X6w775;
wire E7w775, L7w775, S7w775, Z7w775, G8w775, N8w775, U8w775, B9w775, I9w775, P9w775;
wire W9w775, Daw775, Kaw775, Raw775, Yaw775, Fbw775, Mbw775, Tbw775, Acw775, Hcw775;
wire Ocw775, Vcw775, Cdw775, Jdw775, Qdw775, Xdw775, Eew775, Lew775, Sew775, Zew775;
wire Gfw775, Nfw775, Ufw775, Bgw775, Igw775, Pgw775, Wgw775, Dhw775, Khw775, Rhw775;
wire Yhw775, Fiw775, Miw775, Tiw775, Ajw775, Hjw775, Ojw775, Vjw775, Ckw775, Jkw775;
wire Qkw775, Xkw775, Elw775, Llw775, Slw775, Zlw775, Gmw775, Nmw775, Umw775, Bnw775;
wire Inw775, Pnw775, Wnw775, Dow775, Kow775, Row775, Yow775, Fpw775, Mpw775, Tpw775;
wire Aqw775, Hqw775, Oqw775, Vqw775, Crw775, Jrw775, Qrw775, Xrw775, Esw775, Lsw775;
wire Ssw775, Zsw775, Gtw775, Ntw775, Utw775, Buw775, Iuw775, Puw775, Wuw775, Dvw775;
wire Kvw775, Rvw775, Yvw775, Fww775, Mww775, Tww775, Axw775, Hxw775, Oxw775, Vxw775;
wire Cyw775, Jyw775, Qyw775, Xyw775, Ezw775, Lzw775, Szw775, Zzw775, G0x775, N0x775;
wire U0x775, B1x775, I1x775, P1x775, W1x775, D2x775, K2x775, R2x775, Y2x775, F3x775;
wire M3x775, T3x775, A4x775, H4x775, O4x775, V4x775, C5x775, J5x775, Q5x775, X5x775;
wire E6x775, L6x775, S6x775, Z6x775, G7x775, N7x775, U7x775, B8x775, I8x775, P8x775;
wire W8x775, D9x775, K9x775, R9x775, Y9x775, Fax775, Max775, Tax775, Abx775, Hbx775;
wire Obx775, Vbx775, Ccx775, Jcx775, Qcx775, Xcx775, Edx775, Ldx775, Sdx775, Zdx775;
wire Gex775, Nex775, Uex775, Bfx775, Ifx775, Pfx775, Wfx775, Dgx775, Kgx775, Rgx775;
wire Ygx775, Fhx775, Mhx775, Thx775, Aix775, Hix775, Oix775, Vix775, Cjx775, Jjx775;
wire Qjx775, Xjx775, Ekx775, Lkx775, Skx775, Zkx775, Glx775, Nlx775, Ulx775, Bmx775;
wire Imx775, Pmx775, Wmx775, Dnx775, Knx775, Rnx775, Ynx775, Fox775, Mox775, Tox775;
wire Apx775, Hpx775, Opx775, Vpx775, Cqx775, Jqx775, Qqx775, Xqx775, Erx775, Lrx775;
wire Srx775, Zrx775, Gsx775, Nsx775, Usx775, Btx775, Itx775, Ptx775, Wtx775, Dux775;
wire Kux775, Rux775, Yux775, Fvx775, Mvx775, Tvx775, Awx775, Hwx775, Owx775, Vwx775;
wire Cxx775, Jxx775, Qxx775, Xxx775, Eyx775, Lyx775, Syx775, Zyx775, Gzx775, Nzx775;
wire Uzx775, B0y775, I0y775, P0y775, W0y775, D1y775, K1y775, R1y775, Y1y775, F2y775;
wire M2y775, T2y775, A3y775, H3y775, O3y775, V3y775, C4y775, J4y775, Q4y775, X4y775;
wire E5y775, L5y775, S5y775, Z5y775, G6y775, N6y775, U6y775, B7y775, I7y775, P7y775;
wire W7y775, D8y775, K8y775, R8y775, Y8y775, F9y775, M9y775, T9y775, Aay775, Hay775;
wire Oay775, Vay775, Cby775, Jby775, Qby775, Xby775, Ecy775, Lcy775, Scy775, Zcy775;
wire Gdy775, Ndy775, Udy775, Bey775, Iey775, Pey775, Wey775, Dfy775, Kfy775, Rfy775;
wire Yfy775, Fgy775, Mgy775, Tgy775, Ahy775, Hhy775, Ohy775, Vhy775, Ciy775, Jiy775;
wire Qiy775, Xiy775, Ejy775, Ljy775, Sjy775, Zjy775, Gky775, Nky775, Uky775, Bly775;
wire Ily775, Ply775, Wly775, Dmy775, Kmy775, Rmy775, Ymy775, Fny775, Mny775, Tny775;
wire Aoy775, Hoy775, Ooy775, Voy775, Cpy775, Jpy775, Qpy775, Xpy775, Eqy775, Lqy775;
wire Sqy775, Zqy775, Gry775, Nry775, Ury775, Bsy775, Isy775, Psy775, Wsy775, Dty775;
wire Kty775, Rty775, Yty775, Fuy775, Muy775, Tuy775, Avy775, Hvy775, Ovy775, Vvy775;
wire Cwy775, Jwy775, Qwy775, Xwy775, Exy775, Lxy775, Sxy775, Zxy775, Gyy775, Nyy775;
wire Uyy775, Bzy775, Izy775, Pzy775, Wzy775, D0z775, K0z775, R0z775, Y0z775, F1z775;
wire M1z775, T1z775, A2z775, H2z775, O2z775, V2z775, C3z775, J3z775, Q3z775, X3z775;
wire E4z775, L4z775, S4z775, Z4z775, G5z775, N5z775, U5z775, B6z775, I6z775, P6z775;
wire W6z775, D7z775, K7z775, R7z775, Y7z775, F8z775, M8z775, T8z775, A9z775, H9z775;
wire O9z775, V9z775, Caz775, Jaz775, Qaz775, Xaz775, Ebz775, Lbz775, Sbz775, Zbz775;
wire Gcz775, Ncz775, Ucz775, Bdz775, Idz775, Pdz775, Wdz775, Dez775, Kez775, Rez775;
wire Yez775, Ffz775, Mfz775, Tfz775, Agz775, Hgz775, Ogz775, Vgz775, Chz775, Jhz775;
wire Qhz775, Xhz775, Eiz775, Liz775, Siz775, Ziz775, Gjz775, Njz775, Ujz775, Bkz775;
wire Ikz775, Pkz775, Wkz775, Dlz775, Klz775, Rlz775, Ylz775, Fmz775, Mmz775, Tmz775;
wire Anz775, Hnz775, Onz775, Vnz775, Coz775, Joz775, Qoz775, Xoz775, Epz775, Lpz775;
wire Spz775, Zpz775, Gqz775, Nqz775, Uqz775, Brz775, Irz775, Prz775, Wrz775, Dsz775;
wire Ksz775, Rsz775, Ysz775, Ftz775, Mtz775, Ttz775, Auz775, Huz775, Ouz775, Vuz775;
wire Cvz775, Jvz775, Qvz775, Xvz775, Ewz775, Lwz775, Swz775, Zwz775, Gxz775, Nxz775;
wire Uxz775, Byz775, Iyz775, Pyz775, Wyz775, Dzz775, Kzz775, Rzz775, Yzz775, F00875;
wire M00875, T00875, A10875, H10875, O10875, V10875, C20875, J20875, Q20875, X20875;
wire E30875, L30875, S30875, Z30875, G40875, N40875, U40875, B50875, I50875, P50875;
wire W50875, D60875, K60875, R60875, Y60875, F70875, M70875, T70875, A80875, H80875;
wire O80875, V80875, C90875, J90875, Q90875, X90875, Ea0875, La0875, Sa0875, Za0875;
wire Gb0875, Nb0875, Ub0875, Bc0875, Ic0875, Pc0875, Wc0875, Dd0875, Kd0875, Rd0875;
wire Yd0875, Fe0875, Me0875, Te0875, Af0875, Hf0875, Of0875, Vf0875, Cg0875, Jg0875;
wire Qg0875, Xg0875, Eh0875, Lh0875, Sh0875, Zh0875, Gi0875, Ni0875, Ui0875, Bj0875;
wire Ij0875, Pj0875, Wj0875, Dk0875, Kk0875, Rk0875, Yk0875, Fl0875, Ml0875, Tl0875;
wire Am0875, Hm0875, Om0875, Vm0875, Cn0875, Jn0875, Qn0875, Xn0875, Eo0875, Lo0875;
wire So0875, Zo0875, Gp0875, Np0875, Up0875, Bq0875, Iq0875, Pq0875, Wq0875, Dr0875;
wire Kr0875, Rr0875, Yr0875, Fs0875, Ms0875, Ts0875, At0875, Ht0875, Ot0875, Vt0875;
wire Cu0875, Ju0875, Qu0875, Xu0875, Ev0875, Lv0875, Sv0875, Zv0875, Gw0875, Nw0875;
wire Uw0875, Bx0875, Ix0875, Px0875, Wx0875, Dy0875, Ky0875, Ry0875, Yy0875, Fz0875;
wire Mz0875, Tz0875, A01875, H01875, O01875, V01875, C11875, J11875, Q11875, X11875;
wire E21875, L21875, S21875, Z21875, G31875, N31875, U31875, B41875, I41875, P41875;
wire W41875, D51875, K51875, R51875, Y51875, F61875, M61875, T61875, A71875, H71875;
wire O71875, V71875, C81875, J81875, Q81875, X81875, E91875, L91875, S91875, Z91875;
wire Ga1875, Na1875, Ua1875, Bb1875, Ib1875, Pb1875, Wb1875, Dc1875, Kc1875, Rc1875;
wire Yc1875, Fd1875, Md1875, Td1875, Ae1875, He1875, Oe1875, Ve1875, Cf1875, Jf1875;
wire Qf1875, Xf1875, Eg1875, Lg1875, Sg1875, Zg1875, Gh1875, Nh1875, Uh1875, Bi1875;
wire Ii1875, Pi1875, Wi1875, Dj1875, Kj1875, Rj1875, Yj1875, Fk1875, Mk1875, Tk1875;
wire Al1875, Hl1875, Ol1875, Vl1875, Cm1875, Jm1875, Qm1875, Xm1875, En1875, Ln1875;
wire Sn1875, Zn1875, Go1875, No1875, Uo1875, Bp1875, Ip1875, Pp1875, Wp1875, Dq1875;
wire Kq1875, Rq1875, Yq1875, Fr1875, Mr1875, Tr1875, As1875, Hs1875, Os1875, Vs1875;
wire Ct1875, Jt1875, Qt1875, Xt1875, Eu1875, Lu1875, Su1875, Zu1875, Gv1875, Nv1875;
wire Uv1875, Bw1875, Iw1875, Pw1875, Ww1875, Dx1875, Kx1875, Rx1875, Yx1875, Fy1875;
wire My1875, Ty1875, Az1875, Hz1875, Oz1875, Vz1875, C02875, J02875, Q02875, X02875;
wire E12875, L12875, S12875, Z12875, G22875, N22875, U22875, B32875, I32875, P32875;
wire W32875, D42875, K42875, R42875, Y42875, F52875, M52875, T52875, A62875, H62875;
wire O62875, V62875, C72875, J72875, Q72875, X72875, E82875, L82875, S82875, Z82875;
wire G92875, N92875, U92875, Ba2875, Ia2875, Pa2875, Wa2875, Db2875, Kb2875, Rb2875;
wire Yb2875, Fc2875, Mc2875, Tc2875, Ad2875, Hd2875, Od2875, Vd2875, Ce2875, Je2875;
wire Qe2875, Xe2875, Ef2875, Lf2875, Sf2875, Zf2875, Gg2875, Ng2875, Ug2875, Bh2875;
wire Ih2875, Ph2875, Wh2875, Di2875, Ki2875, Ri2875, Yi2875, Fj2875, Mj2875, Tj2875;
wire Ak2875, Hk2875, Ok2875, Vk2875, Cl2875, Jl2875, Ql2875, Xl2875, Em2875, Lm2875;
wire Sm2875, Zm2875, Gn2875, Nn2875, Un2875, Bo2875, Io2875, Po2875, Wo2875, Dp2875;
wire Kp2875, Rp2875, Yp2875, Fq2875, Mq2875, Tq2875, Ar2875, Hr2875, Or2875, Vr2875;
wire Cs2875, Js2875, Qs2875, Xs2875, Et2875, Lt2875, St2875, Zt2875, Gu2875, Nu2875;
wire Uu2875, Bv2875, Iv2875, Pv2875, Wv2875, Dw2875, Kw2875, Rw2875, Yw2875, Fx2875;
wire Mx2875, Tx2875, Ay2875, Hy2875, Oy2875, Vy2875, Cz2875, Jz2875, Qz2875, Xz2875;
wire E03875, L03875, S03875, Z03875, G13875, N13875, U13875, B23875, I23875, P23875;
wire W23875, D33875, K33875, R33875, Y33875, F43875, M43875, T43875, A53875, H53875;
wire O53875, V53875, C63875, J63875, Q63875, X63875, E73875, L73875, S73875, Z73875;
wire G83875, N83875, U83875, B93875, I93875, P93875, W93875, Da3875, Ka3875, Ra3875;
wire Ya3875, Fb3875, Mb3875, Tb3875, Ac3875, Hc3875, Oc3875, Vc3875, Cd3875, Jd3875;
wire Qd3875, Xd3875, Ee3875, Le3875, Se3875, Ze3875, Gf3875, Nf3875, Uf3875, Bg3875;
wire Ig3875, Pg3875, Wg3875, Dh3875, Kh3875, Rh3875, Yh3875, Fi3875, Mi3875, Ti3875;
wire Aj3875, Hj3875, Oj3875, Vj3875, Ck3875, Jk3875, Qk3875, Xk3875, El3875, Ll3875;
wire Sl3875, Zl3875, Gm3875, Nm3875, Um3875, Bn3875, In3875, Pn3875, Wn3875, Do3875;
wire Ko3875, Ro3875, Yo3875, Fp3875, Mp3875, Tp3875, Aq3875, Hq3875, Oq3875, Vq3875;
wire Cr3875, Jr3875, Qr3875, Xr3875, Es3875, Ls3875, Ss3875, Zs3875, Gt3875, Nt3875;
wire Ut3875, Bu3875, Iu3875, Pu3875, Wu3875, Dv3875, Kv3875, Rv3875, Yv3875, Fw3875;
wire Mw3875, Tw3875, Ax3875, Hx3875, Ox3875, Vx3875, Cy3875, Jy3875, Qy3875, Xy3875;
wire Ez3875, Lz3875, Sz3875, Zz3875, G04875, N04875, U04875, B14875, I14875, P14875;
wire W14875, D24875, K24875, R24875, Y24875, F34875, M34875, T34875, A44875, H44875;
wire O44875, V44875, C54875, J54875, Q54875, X54875, E64875, L64875, S64875, Z64875;
wire G74875, N74875, U74875, B84875, I84875, P84875, W84875, D94875, K94875, R94875;
wire Y94875, Fa4875, Ma4875, Ta4875, Ab4875, Hb4875, Ob4875, Vb4875, Cc4875, Jc4875;
wire Qc4875, Xc4875, Ed4875, Ld4875, Sd4875, Zd4875, Ge4875, Ne4875, Ue4875, Bf4875;
wire If4875, Pf4875, Wf4875, Dg4875, Kg4875, Rg4875, Yg4875, Fh4875, Mh4875, Th4875;
wire Ai4875, Hi4875, Oi4875, Vi4875, Cj4875, Jj4875, Qj4875, Xj4875, Ek4875, Lk4875;
wire Sk4875, Zk4875, Gl4875, Nl4875, Ul4875, Bm4875, Im4875, Pm4875, Wm4875, Dn4875;
wire Kn4875, Rn4875, Yn4875, Fo4875, Mo4875, To4875, Ap4875, Hp4875, Op4875, Vp4875;
wire Cq4875, Jq4875, Qq4875, Xq4875, Er4875, Lr4875, Sr4875, Zr4875, Gs4875, Ns4875;
wire Us4875, Bt4875, It4875, Pt4875, Wt4875, Du4875, Ku4875, Ru4875, Yu4875, Fv4875;
wire Mv4875, Tv4875, Aw4875, Hw4875, Ow4875, Vw4875, Cx4875, Jx4875, Qx4875, Xx4875;
wire Ey4875, Ly4875, Sy4875, Zy4875, Gz4875, Nz4875, Uz4875, B05875, I05875, P05875;
wire W05875, D15875, K15875, R15875, Y15875, F25875, M25875, T25875, A35875, H35875;
wire O35875, V35875, C45875, J45875, Q45875, X45875, E55875, L55875, S55875, Z55875;
wire G65875, N65875, U65875, B75875, I75875, P75875, W75875, D85875, K85875, R85875;
wire Y85875, F95875, M95875, T95875, Aa5875, Ha5875, Oa5875, Va5875, Cb5875, Jb5875;
wire Qb5875, Xb5875, Ec5875, Lc5875, Sc5875, Zc5875, Gd5875, Nd5875, Ud5875, Be5875;
wire Ie5875, Pe5875, We5875, Df5875, Kf5875, Rf5875, Yf5875, Fg5875, Mg5875, Tg5875;
wire Ah5875, Hh5875, Oh5875, Vh5875, Ci5875, Ji5875, Qi5875, Xi5875, Ej5875, Lj5875;
wire Sj5875, Zj5875, Gk5875, Nk5875, Uk5875, Bl5875, Il5875, Pl5875, Wl5875, Dm5875;
wire Km5875, Rm5875, Ym5875, Fn5875, Mn5875, Tn5875, Ao5875, Ho5875, Oo5875, Vo5875;
wire Cp5875, Jp5875, Qp5875, Xp5875, Eq5875, Lq5875, Sq5875, Zq5875, Gr5875, Nr5875;
wire Ur5875, Bs5875, Is5875, Ps5875, Ws5875, Dt5875, Kt5875, Rt5875, Yt5875, Fu5875;
wire Mu5875, Tu5875, Av5875, Hv5875, Ov5875, Vv5875, Cw5875, Jw5875, Qw5875, Xw5875;
wire Ex5875, Lx5875, Sx5875, Zx5875, Gy5875, Ny5875, Uy5875, Bz5875, Iz5875, Pz5875;
wire Wz5875, D06875, K06875, R06875, Y06875, F16875, M16875, T16875, A26875, H26875;
wire O26875, V26875, C36875, J36875, Q36875, X36875, E46875, L46875, S46875, Z46875;
wire G56875, N56875, U56875, B66875, I66875, P66875, W66875, D76875, K76875, R76875;
wire Y76875, F86875, M86875, T86875, A96875, H96875, O96875, V96875, Ca6875, Ja6875;
wire Qa6875, Xa6875, Eb6875, Lb6875, Sb6875, Zb6875, Gc6875, Nc6875, Uc6875, Bd6875;
wire Id6875, Pd6875, Wd6875, De6875, Ke6875, Re6875, Ye6875, Ff6875, Mf6875, Tf6875;
wire Ag6875, Hg6875, Og6875, Vg6875, Ch6875, Jh6875, Qh6875, Xh6875, Ei6875, Li6875;
wire Si6875, Zi6875, Gj6875, Nj6875, Uj6875, Bk6875, Ik6875, Pk6875, Wk6875, Dl6875;
wire Kl6875, Rl6875, Yl6875, Fm6875, Mm6875, Tm6875, An6875, Hn6875, On6875, Vn6875;
wire Co6875, Jo6875, Qo6875, Xo6875, Ep6875, Lp6875, Sp6875, Zp6875, Gq6875, Nq6875;
wire Uq6875, Br6875, Ir6875, Pr6875, Wr6875, Ds6875, Ks6875, Rs6875, Ys6875, Ft6875;
wire Mt6875, Tt6875, Au6875, Hu6875, Ou6875, Vu6875, Cv6875, Jv6875, Qv6875, Xv6875;
wire Ew6875, Lw6875, Sw6875, Zw6875, Gx6875, Nx6875, Ux6875, By6875, Iy6875, Py6875;
wire Wy6875, Dz6875, Kz6875, Rz6875, Yz6875, F07875, M07875, T07875, A17875, H17875;
wire O17875, V17875, C27875, J27875, Q27875, X27875, E37875, L37875, S37875, Z37875;
wire G47875, N47875, U47875, B57875, I57875, P57875, W57875, D67875, K67875, R67875;
wire Y67875, F77875, M77875, T77875, A87875, H87875, O87875, V87875, C97875, J97875;
wire Q97875, X97875, Ea7875, La7875, Sa7875, Za7875, Gb7875, Nb7875, Ub7875, Bc7875;
wire Ic7875, Pc7875, Wc7875, Dd7875, Kd7875, Rd7875, Yd7875, Fe7875, Me7875, Te7875;
wire Af7875, Hf7875, Of7875, Vf7875, Cg7875, Jg7875, Qg7875, Xg7875, Eh7875, Lh7875;
wire Sh7875, Zh7875, Gi7875, Ni7875, Ui7875, Bj7875, Ij7875, Pj7875, Wj7875, Dk7875;
wire Kk7875, Rk7875, Yk7875, Fl7875, Ml7875, Tl7875, Am7875, Hm7875, Om7875, Vm7875;
wire Cn7875, Jn7875, Qn7875, Xn7875, Eo7875, Lo7875, So7875, Zo7875, Gp7875, Np7875;
wire Up7875, Bq7875, Iq7875, Pq7875, Wq7875, Dr7875, Kr7875, Rr7875, Yr7875, Fs7875;
wire Ms7875, Ts7875, At7875, Ht7875, Ot7875, Vt7875, Cu7875, Ju7875, Qu7875, Xu7875;
wire Ev7875, Lv7875, Sv7875, Zv7875, Gw7875, Nw7875, Uw7875, Bx7875, Ix7875, Px7875;
wire Wx7875, Dy7875, Ky7875, Ry7875, Yy7875, Fz7875, Mz7875, Tz7875, A08875, H08875;
wire O08875, V08875, C18875, J18875, Q18875, X18875, E28875, L28875, S28875, Z28875;
wire G38875, N38875, U38875, B48875, I48875, P48875, W48875, D58875, K58875, R58875;
wire Y58875, F68875, M68875, T68875, A78875, H78875, O78875, V78875, C88875, J88875;
wire Q88875, X88875, E98875, L98875, S98875, Z98875, Ga8875, Na8875, Ua8875, Bb8875;
wire Ib8875, Pb8875, Wb8875, Dc8875, Kc8875, Rc8875, Yc8875, Fd8875, Md8875, Td8875;
wire Ae8875, He8875, Oe8875, Ve8875, Cf8875, Jf8875, Qf8875, Xf8875, Eg8875, Lg8875;
wire Sg8875, Zg8875, Gh8875, Nh8875, Uh8875, Bi8875, Ii8875, Pi8875, Wi8875, Dj8875;
wire Kj8875, Rj8875, Yj8875, Fk8875, Mk8875, Tk8875, Al8875, Hl8875, Ol8875, Vl8875;
wire Cm8875, Jm8875, Qm8875, Xm8875, En8875, Ln8875, Sn8875, Zn8875, Go8875, No8875;
wire Uo8875, Bp8875, Ip8875, Pp8875, Wp8875, Dq8875, Kq8875, Rq8875, Yq8875, Fr8875;
wire Mr8875, Tr8875, As8875, Hs8875, Os8875, Vs8875, Ct8875, Jt8875, Qt8875, Xt8875;
wire Eu8875, Lu8875, Su8875, Zu8875, Gv8875, Nv8875, Uv8875, Bw8875, Iw8875, Pw8875;
wire Ww8875, Dx8875, Kx8875, Rx8875, Yx8875, Fy8875, My8875, Ty8875, Az8875, Hz8875;
wire Oz8875, Vz8875, C09875, J09875, Q09875, X09875, E19875, L19875, S19875, Z19875;
wire G29875, N29875, U29875, B39875, I39875, P39875, W39875, D49875, K49875, R49875;
wire Y49875, F59875, M59875, T59875, A69875, H69875, O69875, V69875, C79875, J79875;
wire Q79875, X79875, E89875, L89875, S89875, Z89875, G99875, N99875, U99875, Ba9875;
wire Ia9875, Pa9875, Wa9875, Db9875, Kb9875, Rb9875, Yb9875, Fc9875, Mc9875, Tc9875;
wire Ad9875, Hd9875, Od9875, Vd9875, Ce9875, Je9875, Qe9875, Xe9875, Ef9875, Lf9875;
wire Sf9875, Zf9875, Gg9875, Ng9875, Ug9875, Bh9875, Ih9875, Ph9875, Wh9875, Di9875;
wire Ki9875, Ri9875, Yi9875, Fj9875, Mj9875, Tj9875, Ak9875, Hk9875, Ok9875, Vk9875;
wire Cl9875, Jl9875, Ql9875, Xl9875, Em9875, Lm9875, Sm9875, Zm9875, Gn9875, Nn9875;
wire Un9875, Bo9875, Io9875, Po9875, Wo9875, Dp9875, Kp9875, Rp9875, Yp9875, Fq9875;
wire Mq9875, Tq9875, Ar9875, Hr9875, Or9875, Vr9875, Cs9875, Js9875, Qs9875, Xs9875;
wire Et9875, Lt9875, St9875, Zt9875, Gu9875, Nu9875, Uu9875, Bv9875, Iv9875, Pv9875;
wire Wv9875, Dw9875, Kw9875, Rw9875, Yw9875, Fx9875, Mx9875, Tx9875, Ay9875, Hy9875;
wire Oy9875, Vy9875, Cz9875, Jz9875, Qz9875, Xz9875, E0a875, L0a875, S0a875, Z0a875;
wire G1a875, N1a875, U1a875, B2a875, I2a875, P2a875, W2a875, D3a875, K3a875, R3a875;
wire Y3a875, F4a875, M4a875, T4a875, A5a875, H5a875, O5a875, V5a875, C6a875, J6a875;
wire Q6a875, X6a875, E7a875, L7a875, S7a875, Z7a875, G8a875, N8a875, U8a875, B9a875;
wire I9a875, P9a875, W9a875, Daa875, Kaa875, Raa875, Yaa875, Fba875, Mba875, Tba875;
wire Aca875, Hca875, Oca875, Vca875, Cda875, Jda875, Qda875, Xda875, Eea875, Lea875;
wire Sea875, Zea875, Gfa875, Nfa875, Ufa875, Bga875, Iga875, Pga875, Wga875, Dha875;
wire Kha875, Rha875, Yha875, Fia875, Mia875, Tia875, Aja875, Hja875, Oja875, Vja875;
wire Cka875, Jka875, Qka875, Xka875, Ela875, Lla875, Sla875, Zla875, Gma875, Nma875;
wire Uma875, Bna875, Ina875, Pna875, Wna875, Doa875, Koa875, Roa875, Yoa875, Fpa875;
wire Mpa875, Tpa875, Aqa875, Hqa875, Oqa875, Vqa875, Cra875, Jra875, Qra875, Xra875;
wire Esa875, Lsa875, Ssa875, Zsa875, Gta875, Nta875, Uta875, Bua875, Iua875, Pua875;
wire Wua875, Dva875, Kva875, Rva875, Yva875, Fwa875, Mwa875, Twa875, Axa875, Hxa875;
wire Oxa875, Vxa875, Cya875, Jya875, Qya875, Xya875, Eza875, Lza875, Sza875, Zza875;
wire G0b875, N0b875, U0b875, B1b875, I1b875, P1b875, W1b875, D2b875, K2b875, R2b875;
wire Y2b875, F3b875, M3b875, T3b875, A4b875, H4b875, O4b875, V4b875, C5b875, J5b875;
wire Q5b875, X5b875, E6b875, L6b875, S6b875, Z6b875, G7b875, N7b875, U7b875, B8b875;
wire I8b875, P8b875, W8b875, D9b875, K9b875, R9b875, Y9b875, Fab875, Mab875, Tab875;
wire Abb875, Hbb875, Obb875, Vbb875, Ccb875, Jcb875, Qcb875, Xcb875, Edb875, Ldb875;
wire Sdb875, Zdb875, Geb875, Neb875, Ueb875, Bfb875, Ifb875, Pfb875, Wfb875, Dgb875;
wire Kgb875, Rgb875, Ygb875, Fhb875, Mhb875, Thb875, Aib875, Hib875, Oib875, Vib875;
wire Cjb875, Jjb875, Qjb875, Xjb875, Ekb875, Lkb875, Skb875, Zkb875, Glb875, Nlb875;
wire Ulb875, Bmb875, Imb875, Pmb875, Wmb875, Dnb875, Knb875, Rnb875, Ynb875, Fob875;
wire Mob875, Tob875, Apb875, Hpb875, Opb875, Vpb875, Cqb875, Jqb875, Qqb875, Xqb875;
wire Erb875, Lrb875, Srb875, Zrb875, Gsb875, Nsb875, Usb875, Btb875, Itb875, Ptb875;
wire Wtb875, Dub875, Kub875, Rub875, Yub875, Fvb875, Mvb875, Tvb875, Awb875, Hwb875;
wire Owb875, Vwb875, Cxb875, Jxb875, Qxb875, Xxb875, Eyb875, Lyb875, Syb875, Zyb875;
wire Gzb875, Nzb875, Uzb875, B0c875, I0c875, P0c875, W0c875, D1c875, K1c875, R1c875;
wire Y1c875, F2c875, M2c875, T2c875, A3c875, H3c875, O3c875, V3c875, C4c875, J4c875;
wire Q4c875, X4c875, E5c875, L5c875, S5c875, Z5c875, G6c875, N6c875, U6c875, B7c875;
wire I7c875, P7c875, W7c875, D8c875, K8c875, R8c875, Y8c875, F9c875, M9c875, T9c875;
wire Aac875, Hac875, Oac875, Vac875, Cbc875, Jbc875, Qbc875, Xbc875, Ecc875, Lcc875;
wire Scc875, Zcc875, Gdc875, Ndc875, Udc875, Bec875, Iec875, Pec875, Wec875, Dfc875;
wire Kfc875, Rfc875, Yfc875, Fgc875, Mgc875, Tgc875, Ahc875, Hhc875, Ohc875, Vhc875;
wire Cic875, Jic875, Qic875, Xic875, Ejc875, Ljc875, Sjc875, Zjc875, Gkc875, Nkc875;
wire Ukc875, Blc875, Ilc875, Plc875, Wlc875, Dmc875, Kmc875, Rmc875, Ymc875, Fnc875;
wire Mnc875, Tnc875, Aoc875, Hoc875, Ooc875, Voc875, Cpc875, Jpc875, Qpc875, Xpc875;
wire Eqc875, Lqc875, Sqc875, Zqc875, Grc875, Nrc875, Urc875, Bsc875, Isc875, Psc875;
wire Wsc875, Dtc875, Ktc875, Rtc875, Ytc875, Fuc875, Muc875, Tuc875, Avc875, Hvc875;
wire Ovc875, Vvc875, Cwc875, Jwc875, Qwc875, Xwc875, Exc875, Lxc875, Sxc875, Zxc875;
wire Gyc875, Nyc875, Uyc875, Bzc875, Izc875, Pzc875, Wzc875, D0d875, K0d875, R0d875;
wire Y0d875, F1d875, M1d875, T1d875, A2d875, H2d875, O2d875, V2d875, C3d875, J3d875;
wire Q3d875, X3d875, E4d875, L4d875, S4d875, Z4d875, G5d875, N5d875, U5d875, B6d875;
wire I6d875, P6d875, W6d875, D7d875, K7d875, R7d875, Y7d875, F8d875, M8d875, T8d875;
wire A9d875, H9d875, O9d875, V9d875, Cad875, Jad875, Qad875, Xad875, Ebd875, Lbd875;
wire Sbd875, Zbd875, Gcd875, Ncd875, Ucd875, Bdd875, Idd875, Pdd875, Wdd875, Ded875;
wire Ked875, Red875, Yed875, Ffd875, Mfd875, Tfd875, Agd875, Hgd875, Ogd875, Vgd875;
wire Chd875, Jhd875, Qhd875, Xhd875, Eid875, Lid875, Sid875, Zid875, Gjd875, Njd875;
wire Ujd875, Bkd875, Ikd875, Pkd875, Wkd875, Dld875, Kld875, Rld875, Yld875, Fmd875;
wire Mmd875, Tmd875, And875, Hnd875, Ond875, Vnd875, Cod875, Jod875, Qod875, Xod875;
wire Epd875, Lpd875, Spd875, Zpd875, Gqd875, Nqd875, Uqd875, Brd875, Ird875, Prd875;
wire Wrd875, Dsd875, Ksd875, Rsd875, Ysd875, Ftd875, Mtd875, Ttd875, Aud875, Hud875;
wire Oud875, Vud875, Cvd875, Jvd875, Qvd875, Xvd875, Ewd875, Lwd875, Swd875, Zwd875;
wire Gxd875, Nxd875, Uxd875, Byd875, Iyd875, Pyd875, Wyd875, Dzd875, Kzd875, Rzd875;
wire Yzd875, F0e875, M0e875, T0e875, A1e875, H1e875, O1e875, V1e875, C2e875, J2e875;
wire Q2e875, X2e875, E3e875, L3e875, S3e875, Z3e875, G4e875, N4e875, U4e875, B5e875;
wire I5e875, P5e875, W5e875, D6e875, K6e875, R6e875, Y6e875, F7e875, M7e875, T7e875;
wire A8e875, H8e875, O8e875, V8e875, C9e875, J9e875, Q9e875, X9e875, Eae875, Lae875;
wire Sae875, Zae875, Gbe875, Nbe875, Ube875, Bce875, Ice875, Pce875, Wce875, Dde875;
wire Kde875, Rde875, Yde875, Fee875, Mee875, Tee875, Afe875, Hfe875, Ofe875, Vfe875;
wire Cge875, Jge875, Qge875, Xge875, Ehe875, Lhe875, She875, Zhe875, Gie875, Nie875;
wire Uie875, Bje875, Ije875, Pje875, Wje875, Dke875, Kke875, Rke875, Yke875, Fle875;
wire Mle875, Tle875, Ame875, Hme875, Ome875, Vme875, Cne875, Jne875, Qne875, Xne875;
wire Eoe875, Loe875, Soe875, Zoe875, Gpe875, Npe875, Upe875, Bqe875, Iqe875, Pqe875;
wire Wqe875, Dre875, Kre875, Rre875, Yre875, Fse875, Mse875, Tse875, Ate875, Hte875;
wire Ote875, Vte875, Cue875, Jue875, Que875, Xue875, Eve875, Lve875, Sve875, Zve875;
wire Gwe875, Nwe875, Uwe875, Bxe875, Ixe875, Pxe875, Wxe875, Dye875, Kye875, Rye875;
wire Yye875, Fze875, Mze875, Tze875, A0f875, H0f875, O0f875, V0f875, C1f875, J1f875;
wire Q1f875, X1f875, E2f875, L2f875, S2f875, Z2f875, G3f875, N3f875, U3f875, B4f875;
wire I4f875, Ycgk85, Fdgk85, Mdgk85, Tdgk85, Aegk85, Hegk85, Oegk85, Vegk85, Cfgk85;
wire Jfgk85, Qfgk85, Xfgk85, Eggk85, Lggk85, Sggk85, Zggk85, Ghgk85, Nhgk85, Uhgk85;
wire Bigk85, Iigk85, Pigk85, Wigk85, Djgk85, Kjgk85, Rjgk85, Yjgk85, Fkgk85, Mkgk85;
wire Tkgk85, Algk85, Hlgk85, Olgk85, Vlgk85, Cmgk85, Jmgk85, Qmgk85, Xmgk85, Engk85;
wire Lngk85, Sngk85, Zngk85, Gogk85, Nogk85, Uogk85, Bpgk85, Ipgk85, Ppgk85, Wpgk85;
wire Dqgk85, Kqgk85, Rqgk85, Yqgk85, Frgk85, Mrgk85, Trgk85, Asgk85, Hsgk85, Osgk85;
wire Vsgk85, Ctgk85, Jtgk85, Qtgk85, Xtgk85, Eugk85, Lugk85, Sugk85, Zugk85, Gvgk85;
wire Nvgk85, Uvgk85, Bwgk85, Iwgk85, Pwgk85, Wwgk85, Dxgk85, Kxgk85, Rxgk85, Yxgk85;
wire Fygk85, Mygk85, Tygk85, Azgk85, Hzgk85, Ozgk85, Vzgk85, C0hk85, J0hk85, Q0hk85;
wire X0hk85, E1hk85, L1hk85, S1hk85, Z1hk85, G2hk85, N2hk85, U2hk85, B3hk85, I3hk85;
wire P3hk85, W3hk85, D4hk85, K4hk85, R4hk85, Y4hk85, F5hk85, M5hk85, T5hk85, A6hk85;
wire H6hk85, O6hk85, V6hk85, C7hk85, J7hk85, Q7hk85, X7hk85, E8hk85, L8hk85, S8hk85;
wire Z8hk85, G9hk85, N9hk85, U9hk85, Bahk85, Iahk85, Pahk85, Wahk85, Dbhk85, Kbhk85;
wire Rbhk85, Ybhk85, Fchk85, Mchk85, Tchk85, Adhk85, Hdhk85, Odhk85, Vdhk85, Cehk85;
wire Jehk85, Qehk85, Xehk85, Efhk85, Lfhk85, Sfhk85, Zfhk85, Gghk85, Nghk85, Ughk85;
wire Bhhk85, Ihhk85, Phhk85, Whhk85, Dihk85, Kihk85, Rihk85, Yihk85, Fjhk85, Mjhk85;
wire Tjhk85, Akhk85, Hkhk85, Okhk85, Vkhk85, Clhk85, Jlhk85, Qlhk85, Xlhk85, Emhk85;
wire Lmhk85, Smhk85, Zmhk85, Gnhk85, Nnhk85, Unhk85, Bohk85, Iohk85, Pohk85, Wohk85;
wire Dphk85, Kphk85, Rphk85, Yphk85, Fqhk85, Mqhk85, Tqhk85, Arhk85, Hrhk85, Orhk85;
wire Vrhk85, Cshk85, Jshk85, Qshk85, Xshk85, Ethk85, Lthk85, Sthk85, Zthk85, Guhk85;
wire Nuhk85, Uuhk85, Bvhk85, Ivhk85, Pvhk85, Wvhk85, Dwhk85, Kwhk85, Rwhk85, Ywhk85;
wire Fxhk85, Mxhk85, Txhk85, Ayhk85, Hyhk85, Oyhk85, Vyhk85, Czhk85, Jzhk85, Qzhk85;
wire Xzhk85, E0ik85, L0ik85, S0ik85, Z0ik85, G1ik85, N1ik85, U1ik85, B2ik85, I2ik85;
wire P2ik85, W2ik85, D3ik85, K3ik85, R3ik85, Y3ik85, F4ik85, M4ik85, T4ik85, A5ik85;
wire H5ik85, O5ik85, V5ik85, C6ik85, J6ik85, Q6ik85, X6ik85, E7ik85, L7ik85, S7ik85;
wire Z7ik85, G8ik85, N8ik85, U8ik85, B9ik85, I9ik85, P9ik85, W9ik85, Daik85, Kaik85;
wire Raik85, Yaik85, Fbik85, Mbik85, Tbik85, Acik85, Hcik85, Ocik85, Vcik85, Cdik85;
wire Jdik85, Qdik85, Xdik85, Eeik85, Leik85, Seik85, Zeik85, Gfik85, Nfik85, Ufik85;
wire Bgik85, Igik85, Pgik85, Wgik85, Dhik85, Khik85, Rhik85, Yhik85, Fiik85, Miik85;
wire Tiik85, Ajik85, Hjik85, Ojik85, Vjik85, Ckik85, Jkik85, Qkik85, Xkik85, Elik85;
wire Llik85, Slik85, Zlik85, Gmik85, Nmik85, Umik85, Bnik85, Inik85, Pnik85, Wnik85;
wire Doik85, Koik85, Roik85, Yoik85, Fpik85, Mpik85, Tpik85, Aqik85, Hqik85, Oqik85;
wire Vqik85, Crik85, Jrik85, Qrik85, Xrik85, Esik85, Lsik85, Ssik85, Zsik85, Gtik85;
wire Ntik85, Utik85, Buik85, Iuik85, Puik85, Wuik85, Dvik85, Kvik85, Rvik85, Yvik85;
wire Fwik85, Mwik85, Twik85, Axik85, Hxik85, Oxik85, Vxik85, Cyik85, Jyik85, Qyik85;
wire Xyik85, Ezik85, Lzik85, Szik85, Zzik85, G0jk85, N0jk85, U0jk85, B1jk85, I1jk85;
wire P1jk85, W1jk85, D2jk85, K2jk85, R2jk85, Y2jk85, F3jk85, M3jk85, T3jk85, A4jk85;
wire H4jk85, O4jk85, V4jk85, C5jk85, J5jk85, Q5jk85, X5jk85, E6jk85, L6jk85, S6jk85;
wire Z6jk85, G7jk85, N7jk85, U7jk85, B8jk85, I8jk85, P8jk85, W8jk85, D9jk85, K9jk85;
wire R9jk85, Y9jk85, Fajk85, Majk85, Tajk85, Abjk85, Hbjk85, Objk85, Vbjk85, Ccjk85;
wire Jcjk85, Qcjk85, Xcjk85, Edjk85, Ldjk85, Sdjk85, Zdjk85, Gejk85, Nejk85, Uejk85;
wire Bfjk85, Ifjk85, Pfjk85, Wfjk85, Dgjk85, Kgjk85, Rgjk85, Ygjk85, Fhjk85, Mhjk85;
wire Thjk85, Aijk85, Hijk85, Oijk85, Vijk85, Cjjk85, Jjjk85, Qjjk85, Xjjk85, Ekjk85;
wire Lkjk85, Skjk85, Zkjk85, Gljk85, Nljk85, Uljk85, Bmjk85, Imjk85, Pmjk85, Wmjk85;
wire Dnjk85, Knjk85, Rnjk85, Ynjk85, Fojk85, Mojk85, Tojk85, Apjk85, Hpjk85, Opjk85;
wire Vpjk85, Cqjk85, Jqjk85, Qqjk85, Xqjk85, Erjk85, Lrjk85, Srjk85, Zrjk85, Gsjk85;
wire Nsjk85, Usjk85, Btjk85, Itjk85, Ptjk85, Wtjk85, Dujk85, Kujk85, Rujk85, Yujk85;
wire Fvjk85, Mvjk85, Tvjk85, Awjk85, Hwjk85, Owjk85, Vwjk85, Cxjk85, Jxjk85, Qxjk85;
wire Xxjk85, Eyjk85, Lyjk85, Syjk85, Zyjk85, Gzjk85, Nzjk85, Uzjk85, B0kk85, I0kk85;
wire P0kk85, W0kk85, D1kk85, K1kk85, R1kk85, Y1kk85, F2kk85, M2kk85, T2kk85, A3kk85;
wire H3kk85, O3kk85, V3kk85, C4kk85, J4kk85, Q4kk85, X4kk85, E5kk85, L5kk85, S5kk85;
wire Z5kk85, G6kk85, N6kk85, U6kk85, B7kk85, I7kk85, P7kk85, W7kk85, D8kk85, K8kk85;
wire R8kk85, Y8kk85, F9kk85, M9kk85, T9kk85, Aakk85, Hakk85, Oakk85, Vakk85, Cbkk85;
wire Jbkk85, Qbkk85, Xbkk85, Eckk85, Lckk85, Sckk85, Zckk85, Gdkk85, Ndkk85, Udkk85;
wire Bekk85, Iekk85, Pekk85, Wekk85, Dfkk85, Kfkk85, Rfkk85, Yfkk85, Fgkk85, Mgkk85;
wire Tgkk85, Ahkk85, Hhkk85, Ohkk85, Vhkk85, Cikk85, Jikk85, Qikk85, Xikk85, Ejkk85;
wire Ljkk85, Sjkk85, Zjkk85, Gkkk85, Nkkk85, Ukkk85, Blkk85, Ilkk85, Plkk85, Wlkk85;
wire Dmkk85, Kmkk85, Rmkk85, Ymkk85, Fnkk85, Mnkk85, Tnkk85, Aokk85, Hokk85, Ookk85;
wire Vokk85, Cpkk85, Jpkk85, Qpkk85, Xpkk85, Eqkk85, Lqkk85, Sqkk85, Zqkk85, Grkk85;
wire Nrkk85, Urkk85, Bskk85, Iskk85, Pskk85, Wskk85, Dtkk85, Ktkk85, Rtkk85, Ytkk85;
wire Fukk85, Mukk85, Tukk85, Avkk85, Hvkk85, Ovkk85, Vvkk85, Cwkk85, Jwkk85, Qwkk85;
wire Xwkk85, Exkk85, Lxkk85, Sxkk85, Zxkk85, Gykk85, Nykk85, Uykk85, Bzkk85, Izkk85;
wire Pzkk85, Wzkk85, D0lk85, K0lk85, R0lk85, Y0lk85, F1lk85, M1lk85, T1lk85, A2lk85;
wire H2lk85, O2lk85, V2lk85, C3lk85, J3lk85, Q3lk85, X3lk85, E4lk85, L4lk85, S4lk85;
wire Z4lk85, G5lk85, N5lk85, U5lk85, B6lk85, I6lk85, P6lk85, W6lk85, D7lk85, K7lk85;
wire R7lk85, Y7lk85, F8lk85, M8lk85, T8lk85, A9lk85, H9lk85, O9lk85, V9lk85, Calk85;
wire Jalk85, Qalk85, Xalk85, Eblk85, Lblk85, Sblk85, Zblk85, Gclk85, Nclk85, Uclk85;
wire Bdlk85, Idlk85, Pdlk85, Wdlk85, Delk85, Kelk85, Relk85, Yelk85, Fflk85, Mflk85;
wire Tflk85, Aglk85, Hglk85, Oglk85, Vglk85, Chlk85, Jhlk85, Qhlk85, Xhlk85, Eilk85;
wire Lilk85, Silk85, Zilk85, Gjlk85, Njlk85, Ujlk85, Bklk85, Iklk85, Pklk85, Wklk85;
wire Dllk85, Kllk85, Rllk85, Yllk85, Fmlk85, Mmlk85, Tmlk85, Anlk85, Hnlk85, Onlk85;
wire Vnlk85, Colk85, Jolk85, Qolk85, Xolk85, Eplk85, Lplk85, Splk85, Zplk85, Gqlk85;
wire Nqlk85, Uqlk85, Brlk85, Irlk85, Prlk85, Wrlk85, Dslk85, Kslk85, Rslk85, Yslk85;
wire Ftlk85, Mtlk85, Ttlk85, Aulk85, Hulk85, Oulk85, Vulk85, Cvlk85, Jvlk85, Qvlk85;
wire Xvlk85, Ewlk85, Lwlk85, Swlk85, Zwlk85, Gxlk85, Nxlk85, Uxlk85, Bylk85, Iylk85;
wire Pylk85, Wylk85, Dzlk85, Kzlk85, Rzlk85, Yzlk85, F0mk85, M0mk85, T0mk85, A1mk85;
wire H1mk85, O1mk85, V1mk85, C2mk85, J2mk85, Q2mk85, X2mk85, E3mk85, L3mk85, S3mk85;
wire Z3mk85, G4mk85, N4mk85, U4mk85, B5mk85, I5mk85, P5mk85, W5mk85, D6mk85, K6mk85;
wire R6mk85, Y6mk85, F7mk85, M7mk85, T7mk85, A8mk85, H8mk85, O8mk85, V8mk85, C9mk85;
wire J9mk85, Q9mk85, X9mk85, Eamk85, Lamk85, Samk85, Zamk85, Gbmk85, Nbmk85, Ubmk85;
wire Bcmk85, Icmk85, Pcmk85, Wcmk85, Ddmk85, Kdmk85, Rdmk85, Ydmk85, Femk85, Memk85;
wire Temk85, Afmk85, Hfmk85, Ofmk85, Vfmk85, Cgmk85, Jgmk85, Qgmk85, Xgmk85, Ehmk85;
wire Lhmk85, Shmk85, Zhmk85, Gimk85, Nimk85, Uimk85, Bjmk85, Ijmk85, Pjmk85, Wjmk85;
wire Dkmk85, Kkmk85, Rkmk85, Ykmk85, Flmk85, Mlmk85, Tlmk85, Ammk85, Hmmk85, Ommk85;
wire Vmmk85, Cnmk85, Jnmk85, Qnmk85, Xnmk85, Eomk85, Lomk85, Somk85, Zomk85, Gpmk85;
wire Npmk85, Upmk85, Bqmk85, Iqmk85, Pqmk85, Wqmk85, Drmk85, Krmk85, Rrmk85, Yrmk85;
wire Fsmk85, Msmk85, Tsmk85, Atmk85, Htmk85, Otmk85, Vtmk85, Cumk85, Jumk85, Qumk85;
wire Xumk85, Evmk85, Lvmk85, Svmk85, Zvmk85, Gwmk85, Nwmk85, Uwmk85, Bxmk85, Ixmk85;
wire Pxmk85, Wxmk85, Dymk85, Kymk85, Rymk85, Yymk85, Fzmk85, Mzmk85, Tzmk85, A0nk85;
wire H0nk85, O0nk85, V0nk85, C1nk85, J1nk85, Q1nk85, X1nk85, E2nk85, L2nk85, S2nk85;
wire Z2nk85, G3nk85, N3nk85, U3nk85, B4nk85, I4nk85, P4nk85, W4nk85, D5nk85, K5nk85;
wire R5nk85, Y5nk85, F6nk85, M6nk85, T6nk85, A7nk85, H7nk85, O7nk85, V7nk85, C8nk85;
wire J8nk85, Q8nk85, X8nk85, E9nk85, L9nk85, S9nk85, Z9nk85, Gank85, Nank85, Uank85;
wire Bbnk85, Ibnk85, Pbnk85, Wbnk85, Dcnk85, Kcnk85, Rcnk85, Ycnk85, Fdnk85, Mdnk85;
wire Tdnk85, Aenk85, Henk85, Oenk85, Venk85, Cfnk85, Jfnk85, Qfnk85, Xfnk85, Egnk85;
wire Lgnk85, Sgnk85, Zgnk85, Ghnk85, Nhnk85, Uhnk85, Bink85, Iink85, Pink85, Wink85;
wire Djnk85, Kjnk85, Rjnk85, Yjnk85, Fknk85, Mknk85, Tknk85, Alnk85, Hlnk85, Olnk85;
wire Vlnk85, Cmnk85, Jmnk85, Qmnk85, Xmnk85, Ennk85, Lnnk85, Snnk85, Znnk85, Gonk85;
wire Nonk85, Uonk85, Bpnk85, Ipnk85, Ppnk85, Wpnk85, Dqnk85, Kqnk85, Rqnk85, Yqnk85;
wire Frnk85, Mrnk85, Trnk85, Asnk85, Hsnk85, Osnk85, Vsnk85, Ctnk85, Jtnk85, Qtnk85;
wire Xtnk85, Eunk85, Lunk85, Sunk85, Zunk85, Gvnk85, Nvnk85, Uvnk85, Bwnk85, Iwnk85;
wire Pwnk85, Wwnk85, Dxnk85, Kxnk85, Rxnk85, Yxnk85, Fynk85, Mynk85, Tynk85, Aznk85;
wire Hznk85, Oznk85, Vznk85, C0ok85, J0ok85, Q0ok85, X0ok85, E1ok85, L1ok85, S1ok85;
wire Z1ok85, G2ok85, N2ok85, U2ok85, B3ok85, I3ok85, P3ok85, W3ok85, D4ok85, K4ok85;
wire R4ok85, Y4ok85, F5ok85, M5ok85, T5ok85, A6ok85, H6ok85, O6ok85, V6ok85, C7ok85;
wire J7ok85, Q7ok85, X7ok85, E8ok85, L8ok85, S8ok85, Z8ok85, G9ok85, N9ok85, U9ok85;
wire Baok85, Iaok85, Paok85, Waok85, Dbok85, Kbok85, Rbok85, Ybok85, Fcok85, Mcok85;
wire Tcok85, Adok85, Hdok85, Odok85, Vdok85, Ceok85, Jeok85, Qeok85, Xeok85, Efok85;
wire Lfok85, Sfok85, Zfok85, Ggok85, Ngok85, Ugok85, Bhok85, Ihok85, Phok85, Whok85;
wire Diok85, Kiok85, Riok85, Yiok85, Fjok85, Mjok85, Tjok85, Akok85, Hkok85, Okok85;
wire Vkok85, Clok85, Jlok85, Qlok85, Xlok85, Emok85, Lmok85, Smok85, Zmok85, Gnok85;
wire Nnok85, Unok85, Book85, Iook85, Pook85, Wook85, Dpok85, Kpok85, Rpok85, Ypok85;
wire Fqok85, Mqok85, Tqok85, Arok85, Hrok85, Orok85, Vrok85, Csok85, Jsok85, Qsok85;
wire Xsok85, Etok85, Ltok85, Stok85, Ztok85, Guok85, Nuok85, Uuok85, Bvok85, Ivok85;
wire Pvok85, Wvok85, Dwok85, Kwok85, Rwok85, Ywok85, Fxok85, Mxok85, Txok85, Ayok85;
wire Hyok85, Oyok85, Vyok85, Czok85, Jzok85, Qzok85, Xzok85, E0pk85, L0pk85, S0pk85;
wire Z0pk85, G1pk85, N1pk85, U1pk85, B2pk85, I2pk85, P2pk85, W2pk85, D3pk85, K3pk85;
wire R3pk85, Y3pk85, F4pk85, M4pk85, T4pk85, A5pk85, H5pk85, O5pk85, V5pk85, C6pk85;
wire J6pk85, Q6pk85, X6pk85, E7pk85, L7pk85, S7pk85, Z7pk85, G8pk85, N8pk85, U8pk85;
wire B9pk85, I9pk85, P9pk85, W9pk85, Dapk85, Kapk85, Rapk85, Yapk85, Fbpk85, Mbpk85;
wire Tbpk85, Acpk85, Hcpk85, Ocpk85, Vcpk85, Cdpk85, Jdpk85, Qdpk85, Xdpk85, Eepk85;
wire Lepk85, Sepk85, Zepk85, Gfpk85, Nfpk85, Ufpk85, Bgpk85, Igpk85, Pgpk85, Wgpk85;
wire Dhpk85, Khpk85, Rhpk85, Yhpk85, Fipk85, Mipk85, Tipk85, Ajpk85, Hjpk85, Ojpk85;
wire Vjpk85, Ckpk85, Jkpk85, Qkpk85, Xkpk85, Elpk85, Llpk85, Slpk85, Zlpk85, Gmpk85;
wire Nmpk85, Umpk85, Bnpk85, Inpk85, Pnpk85, Wnpk85, Dopk85, Kopk85, Ropk85, Yopk85;
wire Fppk85, Mppk85, Tppk85, Aqpk85, Hqpk85, Oqpk85, Vqpk85, Crpk85, Jrpk85, Qrpk85;
wire Xrpk85, Espk85, Lspk85, Sspk85, Zspk85, Gtpk85, Ntpk85, Utpk85, Bupk85, Iupk85;
wire Pupk85, Wupk85, Dvpk85, Kvpk85, Rvpk85, Yvpk85, Fwpk85, Mwpk85, Twpk85, Axpk85;
wire Hxpk85, Oxpk85, Vxpk85, Cypk85, Jypk85, Qypk85, Xypk85, Ezpk85, Lzpk85, Szpk85;
wire Zzpk85, G0qk85, N0qk85, U0qk85, B1qk85, I1qk85, P1qk85, W1qk85, D2qk85, K2qk85;
wire R2qk85, Y2qk85, F3qk85, M3qk85, T3qk85, A4qk85, H4qk85, O4qk85, V4qk85, C5qk85;
wire J5qk85, Q5qk85, X5qk85, E6qk85, L6qk85, S6qk85, Z6qk85, G7qk85, N7qk85, U7qk85;
wire B8qk85, I8qk85, P8qk85, W8qk85, D9qk85, K9qk85, R9qk85, Y9qk85, Faqk85, Maqk85;
wire Taqk85, Abqk85, Hbqk85, Obqk85, Vbqk85, Ccqk85, Jcqk85, Qcqk85, Xcqk85, Edqk85;
wire Ldqk85, Sdqk85, Zdqk85, Geqk85, Neqk85, Ueqk85, Bfqk85, Ifqk85, Pfqk85, Wfqk85;
wire Dgqk85, Kgqk85, Rgqk85, Ygqk85, Fhqk85, Mhqk85, Thqk85, Aiqk85, Hiqk85, Oiqk85;
wire Viqk85, Cjqk85, Jjqk85, Qjqk85, Xjqk85, Ekqk85, Lkqk85, Skqk85, Zkqk85, Glqk85;
wire Nlqk85, Ulqk85, Bmqk85, Imqk85, Pmqk85, Wmqk85, Dnqk85, Knqk85, Rnqk85, Ynqk85;
wire Foqk85, Moqk85, Toqk85, Apqk85, Hpqk85, Opqk85, Vpqk85, Cqqk85, Jqqk85, Qqqk85;
wire Xqqk85, Erqk85, Lrqk85, Srqk85, Zrqk85, Gsqk85, Nsqk85, Usqk85, Btqk85, Itqk85;
wire Ptqk85, Wtqk85, Duqk85, Kuqk85, Ruqk85, Yuqk85, Fvqk85, Mvqk85, Tvqk85, Awqk85;
wire Hwqk85, Owqk85, Vwqk85, Cxqk85, Jxqk85, Qxqk85, Xxqk85, Eyqk85, Lyqk85, Syqk85;
wire Zyqk85, Gzqk85, Nzqk85, Uzqk85, B0rk85, I0rk85, P0rk85, W0rk85, D1rk85, K1rk85;
wire R1rk85, Y1rk85, F2rk85, M2rk85, T2rk85, A3rk85, H3rk85, O3rk85, V3rk85, C4rk85;
wire J4rk85, Q4rk85, X4rk85, E5rk85, L5rk85, S5rk85, Z5rk85, G6rk85, N6rk85, U6rk85;
wire B7rk85, I7rk85, P7rk85, W7rk85, D8rk85, K8rk85, R8rk85, Y8rk85, F9rk85, M9rk85;
wire T9rk85, Aark85, Hark85, Oark85, Vark85, Cbrk85, Jbrk85, Qbrk85, Xbrk85, Ecrk85;
wire Lcrk85, Scrk85, Zcrk85, Gdrk85, Ndrk85, Udrk85, Berk85, Ierk85, Perk85, Werk85;
wire Dfrk85, Kfrk85, Rfrk85, Yfrk85, Fgrk85, Mgrk85, Tgrk85, Ahrk85, Hhrk85, Ohrk85;
wire Vhrk85, Cirk85, Jirk85, Qirk85, Xirk85, Ejrk85, Ljrk85, Sjrk85, Zjrk85, Gkrk85;
wire Nkrk85, Ukrk85, Blrk85, Ilrk85, Plrk85, Wlrk85, Dmrk85, Kmrk85, Rmrk85, Ymrk85;
wire Fnrk85, Mnrk85, Tnrk85, Aork85, Hork85, Oork85, Vork85, Cprk85, Jprk85, Qprk85;
wire Xprk85, Eqrk85, Lqrk85, Sqrk85, Zqrk85, Grrk85, Nrrk85, Urrk85, Bsrk85, Isrk85;
wire Psrk85, Wsrk85, Dtrk85, Ktrk85, Rtrk85, Ytrk85, Furk85, Murk85, Turk85, Avrk85;
wire Hvrk85, Ovrk85, Vvrk85, Cwrk85, Jwrk85, Qwrk85, Xwrk85, Exrk85, Lxrk85, Sxrk85;
wire Zxrk85, Gyrk85, Nyrk85, Uyrk85, Bzrk85, Izrk85, Pzrk85, Wzrk85, D0sk85, K0sk85;
wire R0sk85, Y0sk85, F1sk85, M1sk85, T1sk85, A2sk85, H2sk85, O2sk85, V2sk85, C3sk85;
wire J3sk85, Q3sk85, X3sk85, E4sk85, L4sk85, S4sk85, Z4sk85, G5sk85, N5sk85, U5sk85;
wire B6sk85, I6sk85, P6sk85, W6sk85, D7sk85, K7sk85, R7sk85, Y7sk85, F8sk85, M8sk85;
wire T8sk85, A9sk85, H9sk85, O9sk85, V9sk85, Cask85, Jask85, Qask85, Xask85, Ebsk85;
wire Lbsk85, Sbsk85, Zbsk85, Gcsk85, Ncsk85, Ucsk85, Bdsk85, Idsk85, Pdsk85, Wdsk85;
wire Desk85, Kesk85, Resk85, Yesk85, Ffsk85, Mfsk85, Tfsk85, Agsk85, Hgsk85, Ogsk85;
wire Vgsk85, Chsk85, Jhsk85, Qhsk85, Xhsk85, Eisk85, Lisk85, Sisk85, Zisk85, Gjsk85;
wire Njsk85, Ujsk85, Bksk85, Iksk85, Pksk85, Wksk85, Dlsk85, Klsk85, Rlsk85, Ylsk85;
wire Fmsk85, Mmsk85, Tmsk85, Ansk85, Hnsk85, Onsk85, Vnsk85, Cosk85, Josk85, Qosk85;
wire Xosk85, Epsk85, Lpsk85, Spsk85, Zpsk85, Gqsk85, Nqsk85, Uqsk85, Brsk85, Irsk85;
wire Prsk85, Wrsk85, Dssk85, Kssk85, Rssk85, Yssk85, Ftsk85, Mtsk85, Ttsk85, Ausk85;
wire Husk85, Ousk85, Vusk85, Cvsk85, Jvsk85, Qvsk85, Xvsk85, Ewsk85, Lwsk85, Swsk85;
wire Zwsk85, Gxsk85, Nxsk85, Uxsk85, Bysk85, Iysk85, Pysk85, Wysk85, Dzsk85, Kzsk85;
wire Rzsk85, Yzsk85, F0tk85, M0tk85, T0tk85, A1tk85, H1tk85, O1tk85, V1tk85, C2tk85;
wire J2tk85, Q2tk85, X2tk85, E3tk85, L3tk85, S3tk85, Z3tk85, G4tk85, N4tk85, U4tk85;
wire B5tk85, I5tk85, P5tk85, W5tk85, D6tk85, K6tk85, R6tk85, Y6tk85, F7tk85, M7tk85;
wire T7tk85, A8tk85, H8tk85, O8tk85, V8tk85, C9tk85, J9tk85, Q9tk85, X9tk85, Eatk85;
wire Latk85, Satk85, Zatk85, Gbtk85, Nbtk85, Ubtk85, Bctk85, Ictk85, Pctk85, Wctk85;
wire Ddtk85, Kdtk85, Rdtk85, Ydtk85, Fetk85, Metk85, Tetk85, Aftk85, Hftk85, Oftk85;
wire Vftk85, Cgtk85, Jgtk85, Qgtk85, Xgtk85, Ehtk85, Lhtk85, Shtk85, Zhtk85, Gitk85;
wire Nitk85, Uitk85, Bjtk85, Ijtk85, Pjtk85, Wjtk85, Dktk85, Kktk85, Rktk85, Yktk85;
wire Fltk85, Mltk85, Tltk85, Amtk85, Hmtk85, Omtk85, Vmtk85, Cntk85, Jntk85, Qntk85;
wire Xntk85, Eotk85, Lotk85, Sotk85, Zotk85, Gptk85, Nptk85, Uptk85, Bqtk85, Iqtk85;
wire Pqtk85, Wqtk85, Drtk85, Krtk85, Rrtk85, Yrtk85, Fstk85, Mstk85, Tstk85, Attk85;
wire Httk85, Ottk85, Vttk85, Cutk85, Jutk85, Qutk85, Xutk85, Evtk85, Lvtk85, Svtk85;
wire Zvtk85, Gwtk85, Nwtk85, Uwtk85, Bxtk85, Ixtk85, Pxtk85, Wxtk85, Dytk85, Kytk85;
wire Rytk85, Yytk85, Fztk85, Mztk85, Tztk85, A0uk85, H0uk85, O0uk85, V0uk85, C1uk85;
wire J1uk85, Q1uk85, X1uk85, E2uk85, L2uk85, S2uk85, Z2uk85, G3uk85, N3uk85, U3uk85;
wire B4uk85, I4uk85, P4uk85, W4uk85, D5uk85, K5uk85, R5uk85, Y5uk85, F6uk85, M6uk85;
wire T6uk85, A7uk85, H7uk85, O7uk85, V7uk85, C8uk85, J8uk85, Q8uk85, X8uk85, E9uk85;
wire L9uk85, S9uk85, Z9uk85, Gauk85, Nauk85, Uauk85, Bbuk85, Ibuk85, Pbuk85, Wbuk85;
wire Dcuk85, Kcuk85, Rcuk85, Ycuk85, Fduk85, Mduk85, Tduk85, Aeuk85, Heuk85, Oeuk85;
wire Veuk85, Cfuk85, Jfuk85, Qfuk85, Xfuk85, Eguk85, Lguk85, Sguk85, Zguk85, Ghuk85;
wire Nhuk85, Uhuk85, Biuk85, Iiuk85, Piuk85, Wiuk85, Djuk85, Kjuk85, Rjuk85, Yjuk85;
wire Fkuk85, Mkuk85, Tkuk85, Aluk85, Hluk85, Oluk85, Vluk85, Cmuk85, Jmuk85, Qmuk85;
wire Xmuk85, Enuk85, Lnuk85, Snuk85, Znuk85, Gouk85, Nouk85, Uouk85, Bpuk85, Ipuk85;
wire Ppuk85, Wpuk85, Dquk85, Kquk85, Rquk85, Yquk85, Fruk85, Mruk85, Truk85, Asuk85;
wire Hsuk85, Osuk85, Vsuk85, Ctuk85, Jtuk85, Qtuk85, Xtuk85, Euuk85, Luuk85, Suuk85;
wire Zuuk85, Gvuk85, Nvuk85, Uvuk85, Bwuk85, Iwuk85, Pwuk85, Wwuk85, Dxuk85, Kxuk85;
wire Rxuk85, Yxuk85, Fyuk85, Myuk85, Tyuk85, Azuk85, Hzuk85, Ozuk85, Vzuk85, C0vk85;
wire J0vk85, Q0vk85, X0vk85, E1vk85, L1vk85, S1vk85, Z1vk85, G2vk85, N2vk85, U2vk85;
wire B3vk85, I3vk85, P3vk85, W3vk85, D4vk85, K4vk85, R4vk85, Y4vk85, F5vk85, M5vk85;
wire T5vk85, A6vk85, H6vk85, O6vk85, V6vk85, C7vk85, J7vk85, Q7vk85, X7vk85, E8vk85;
wire L8vk85, S8vk85, Z8vk85, G9vk85, N9vk85, U9vk85, Bavk85, Iavk85, Pavk85, Wavk85;
wire Dbvk85, Kbvk85, Rbvk85, Ybvk85, Fcvk85, Mcvk85, Tcvk85, Advk85, Hdvk85, Odvk85;
wire Vdvk85, Cevk85, Jevk85, Qevk85, Xevk85, Efvk85, Lfvk85, Sfvk85, Zfvk85, Ggvk85;
wire Ngvk85, Ugvk85, Bhvk85, Ihvk85, Phvk85, Whvk85, Divk85, Kivk85, Rivk85, Yivk85;
wire Fjvk85, Mjvk85, Tjvk85, Akvk85, Hkvk85, Okvk85, Vkvk85, Clvk85, Jlvk85, Qlvk85;
wire Xlvk85, Emvk85, Lmvk85, Smvk85, Zmvk85, Gnvk85, Nnvk85, Unvk85, Bovk85, Iovk85;
wire Povk85, Wovk85, Dpvk85, Kpvk85, Rpvk85, Ypvk85, Fqvk85, Mqvk85, Tqvk85, Arvk85;
wire Hrvk85, Orvk85, Vrvk85, Csvk85, Jsvk85, Qsvk85, Xsvk85, Etvk85, Ltvk85, Stvk85;
wire Ztvk85, Guvk85, Nuvk85, Uuvk85, Bvvk85, Ivvk85, Pvvk85, Wvvk85, Dwvk85, Kwvk85;
wire Rwvk85, Ywvk85, Fxvk85, Mxvk85, Txvk85, Ayvk85, Hyvk85, Oyvk85, Vyvk85, Czvk85;
wire Jzvk85, Qzvk85, Xzvk85, E0wk85, L0wk85, S0wk85, Z0wk85, G1wk85, N1wk85, U1wk85;
wire B2wk85, I2wk85, P2wk85, W2wk85, D3wk85, K3wk85, R3wk85, Y3wk85, F4wk85, M4wk85;
wire T4wk85, A5wk85, H5wk85, O5wk85, V5wk85, C6wk85, J6wk85, Q6wk85, X6wk85, E7wk85;
wire L7wk85, S7wk85, Z7wk85, G8wk85, N8wk85, U8wk85, B9wk85, I9wk85, P9wk85, W9wk85;
wire Dawk85, Kawk85, Rawk85, Yawk85, Fbwk85, Mbwk85, Tbwk85, Acwk85, Hcwk85, Ocwk85;
wire Vcwk85, Cdwk85, Jdwk85, Qdwk85, Xdwk85, Eewk85, Lewk85, Sewk85, Zewk85, Gfwk85;
wire Nfwk85, Ufwk85, Bgwk85, Igwk85, Pgwk85, Wgwk85, Dhwk85, Khwk85, Rhwk85, Yhwk85;
wire Fiwk85, Miwk85, Tiwk85, Ajwk85, Hjwk85, Ojwk85, Vjwk85, Ckwk85, Jkwk85, Qkwk85;
wire Xkwk85, Elwk85, Llwk85, Slwk85, Zlwk85, Gmwk85, Nmwk85, Umwk85, Bnwk85, Inwk85;
wire Pnwk85, Wnwk85, Dowk85, Kowk85, Rowk85, Yowk85, Fpwk85, Mpwk85, Tpwk85, Aqwk85;
wire Hqwk85, Oqwk85, Vqwk85, Crwk85, Jrwk85, Qrwk85, Xrwk85, Eswk85, Lswk85, Sswk85;
wire Zswk85, Gtwk85, Ntwk85, Utwk85, Buwk85, Iuwk85, Puwk85, Wuwk85, Dvwk85, Kvwk85;
wire Rvwk85, Yvwk85, Fwwk85, Mwwk85, Twwk85, Axwk85, Hxwk85, Oxwk85, Vxwk85, Cywk85;
wire Jywk85, Qywk85, Xywk85, Ezwk85, Lzwk85, Szwk85, Zzwk85, G0xk85, N0xk85, U0xk85;
wire B1xk85, I1xk85, P1xk85, W1xk85, D2xk85, K2xk85, R2xk85, Y2xk85, F3xk85, M3xk85;
wire T3xk85, A4xk85, H4xk85, O4xk85, V4xk85, C5xk85, J5xk85, Q5xk85, X5xk85, E6xk85;
wire L6xk85, S6xk85, Z6xk85, G7xk85, N7xk85, U7xk85, B8xk85, I8xk85, P8xk85, W8xk85;
wire D9xk85, K9xk85, R9xk85, Y9xk85, Faxk85, Maxk85, Taxk85, Abxk85, Hbxk85, Obxk85;
wire Vbxk85, Ccxk85, Jcxk85, Qcxk85, Xcxk85, Edxk85, Ldxk85, Sdxk85, Zdxk85, Gexk85;
wire Nexk85, Uexk85, Bfxk85, Ifxk85, Pfxk85, Wfxk85, Dgxk85, Kgxk85, Rgxk85, Ygxk85;
wire Fhxk85, Mhxk85, Thxk85, Aixk85, Hixk85, Oixk85, Vixk85, Cjxk85, Jjxk85, Qjxk85;
wire Xjxk85, Ekxk85, Lkxk85, Skxk85, Zkxk85, Glxk85, Nlxk85, Ulxk85, Bmxk85, Imxk85;
wire Pmxk85, Wmxk85, Dnxk85, Knxk85, Rnxk85, Ynxk85, Foxk85, Moxk85, Toxk85, Apxk85;
wire Hpxk85, Opxk85, Vpxk85, Cqxk85, Jqxk85, Qqxk85, Xqxk85, Erxk85, Lrxk85, Srxk85;
wire Zrxk85, Gsxk85, Nsxk85, Usxk85, Btxk85, Itxk85, Ptxk85, Wtxk85, Duxk85, Kuxk85;
wire Ruxk85, Yuxk85, Fvxk85, Mvxk85, Tvxk85, Awxk85, Hwxk85, Owxk85, Vwxk85, Cxxk85;
wire Jxxk85, Qxxk85, Xxxk85, Eyxk85, Lyxk85, Syxk85, Zyxk85, Gzxk85, Nzxk85, Uzxk85;
wire B0yk85, I0yk85, P0yk85, W0yk85, D1yk85, K1yk85, R1yk85, Y1yk85, F2yk85, M2yk85;
wire T2yk85, A3yk85, H3yk85, O3yk85, V3yk85, C4yk85, J4yk85, Q4yk85, X4yk85, E5yk85;
wire L5yk85, S5yk85, Z5yk85, G6yk85, N6yk85, U6yk85, B7yk85, I7yk85, P7yk85, W7yk85;
wire D8yk85, K8yk85, R8yk85, Y8yk85, F9yk85, M9yk85, T9yk85, Aayk85, Hayk85, Oayk85;
wire Vayk85, Cbyk85, Jbyk85, Qbyk85, Xbyk85, Ecyk85, Lcyk85, Scyk85, Zcyk85, Gdyk85;
wire Ndyk85, Udyk85, Beyk85, Ieyk85, Peyk85, Weyk85, Dfyk85, Kfyk85, Rfyk85, Yfyk85;
wire Fgyk85, Mgyk85, Tgyk85, Ahyk85, Hhyk85, Ohyk85, Vhyk85, Ciyk85, Jiyk85, Qiyk85;
wire Xiyk85, Ejyk85, Ljyk85, Sjyk85, Zjyk85, Gkyk85, Nkyk85, Ukyk85, Blyk85, Ilyk85;
wire Plyk85, Wlyk85, Dmyk85, Kmyk85, Rmyk85, Ymyk85, Fnyk85, Mnyk85, Tnyk85, Aoyk85;
wire Hoyk85, Ooyk85, Voyk85, Cpyk85, Jpyk85, Qpyk85, Xpyk85, Eqyk85, Lqyk85, Sqyk85;
wire Zqyk85, Gryk85, Nryk85, Uryk85, Bsyk85, Isyk85, Psyk85, Wsyk85, Dtyk85, Ktyk85;
wire Rtyk85, Ytyk85, Fuyk85, Muyk85, Tuyk85, Avyk85, Hvyk85, Ovyk85, Vvyk85, Cwyk85;
wire Jwyk85, Qwyk85, Xwyk85, Exyk85, Lxyk85, Sxyk85, Zxyk85, Gyyk85, Nyyk85, Uyyk85;
wire Bzyk85, Izyk85, Pzyk85, Wzyk85, D0zk85, K0zk85, R0zk85, Y0zk85, F1zk85, M1zk85;
wire T1zk85, A2zk85, H2zk85, O2zk85, V2zk85, C3zk85, J3zk85, Q3zk85, X3zk85, E4zk85;
wire L4zk85, S4zk85, Z4zk85, G5zk85, N5zk85, U5zk85, B6zk85, I6zk85, P6zk85, W6zk85;
wire D7zk85, K7zk85, R7zk85, Y7zk85, F8zk85, M8zk85, T8zk85, A9zk85, H9zk85, O9zk85;
wire V9zk85, Cazk85, Jazk85, Qazk85, Xazk85, Ebzk85, Lbzk85, Sbzk85, Zbzk85, Gczk85;
wire Nczk85, Uczk85, Bdzk85, Idzk85, Pdzk85, Wdzk85, Dezk85, Kezk85, Rezk85, Yezk85;
wire Ffzk85, Mfzk85, Tfzk85, Agzk85, Hgzk85, Ogzk85, Vgzk85, Chzk85, Jhzk85, Qhzk85;
wire Xhzk85, Eizk85, Lizk85, Sizk85, Zizk85, Gjzk85, Njzk85, Ujzk85, Bkzk85, Ikzk85;
wire Pkzk85, Wkzk85, Dlzk85, Klzk85, Rlzk85, Ylzk85, Fmzk85, Mmzk85, Tmzk85, Anzk85;
wire Hnzk85, Onzk85, Vnzk85, Cozk85, Jozk85, Qozk85, Xozk85, Epzk85, Lpzk85, Spzk85;
wire Zpzk85, Gqzk85, Nqzk85, Uqzk85, Brzk85, Irzk85, Przk85, Wrzk85, Dszk85, Kszk85;
wire Rszk85, Yszk85, Ftzk85, Mtzk85, Ttzk85, Auzk85, Huzk85, Ouzk85, Vuzk85, Cvzk85;
wire Jvzk85, Qvzk85, Xvzk85, Ewzk85, Lwzk85, Swzk85, Zwzk85, Gxzk85, Nxzk85, Uxzk85;
wire Byzk85, Iyzk85, Pyzk85, Wyzk85, Dzzk85, Kzzk85, Rzzk85, Yzzk85, F00l85, M00l85;
wire T00l85, A10l85, H10l85, O10l85, V10l85, C20l85, J20l85, Q20l85, X20l85, E30l85;
wire L30l85, S30l85, Z30l85, G40l85, N40l85, U40l85, B50l85, I50l85, P50l85, W50l85;
wire D60l85, K60l85, R60l85, Y60l85, F70l85, M70l85, T70l85, A80l85, H80l85, O80l85;
wire V80l85, C90l85, J90l85, Q90l85, X90l85, Ea0l85, La0l85, Sa0l85, Za0l85, Gb0l85;
wire Nb0l85, Ub0l85, Bc0l85, Ic0l85, Pc0l85, Wc0l85, Dd0l85, Kd0l85, Rd0l85, Yd0l85;
wire Fe0l85, Me0l85, Te0l85, Af0l85, Hf0l85, Of0l85, Vf0l85, Cg0l85, Jg0l85, Qg0l85;
wire Xg0l85, Eh0l85, Lh0l85, Sh0l85, Zh0l85, Gi0l85, Ni0l85, Ui0l85, Bj0l85, Ij0l85;
wire Pj0l85, Wj0l85, Dk0l85, Kk0l85, Rk0l85, Yk0l85, Fl0l85, Ml0l85, Tl0l85, Am0l85;
wire Hm0l85, Om0l85, Vm0l85, Cn0l85, Jn0l85, Qn0l85, Xn0l85, Eo0l85, Lo0l85, So0l85;
wire Zo0l85, Gp0l85, Np0l85, Up0l85, Bq0l85, Iq0l85, Pq0l85, Wq0l85, Dr0l85, Kr0l85;
wire Rr0l85, Yr0l85, Fs0l85, Ms0l85, Ts0l85, At0l85, Ht0l85, Ot0l85, Vt0l85, Cu0l85;
wire Ju0l85, Qu0l85, Xu0l85, Ev0l85, Lv0l85, Sv0l85, Zv0l85, Gw0l85, Nw0l85, Uw0l85;
wire Bx0l85, Ix0l85, Px0l85, Wx0l85, Dy0l85, Ky0l85, Ry0l85, Yy0l85, Fz0l85, Mz0l85;
wire Tz0l85, A01l85, H01l85, O01l85, V01l85, C11l85, J11l85, Q11l85, X11l85, E21l85;
wire L21l85, S21l85, Z21l85, G31l85, N31l85, U31l85, B41l85, I41l85, P41l85, W41l85;
wire D51l85, K51l85, R51l85, Y51l85, F61l85, M61l85, T61l85, A71l85, H71l85, O71l85;
wire V71l85, C81l85, J81l85, Q81l85, X81l85, E91l85, L91l85, S91l85, Z91l85, Ga1l85;
wire Na1l85, Ua1l85, Bb1l85, Ib1l85, Pb1l85, Wb1l85, Dc1l85, Kc1l85, Rc1l85, Yc1l85;
wire Fd1l85, Md1l85, Td1l85, Ae1l85, He1l85, Oe1l85, Ve1l85, Cf1l85, Jf1l85, Qf1l85;
wire Xf1l85, Eg1l85, Lg1l85, Sg1l85, Zg1l85, Gh1l85, Nh1l85, Uh1l85, Bi1l85, Ii1l85;
wire Pi1l85, Wi1l85, Dj1l85, Kj1l85, Rj1l85, Yj1l85, Fk1l85, Mk1l85, Tk1l85, Al1l85;
wire Hl1l85, Ol1l85, Vl1l85, Cm1l85, Jm1l85, Qm1l85, Xm1l85, En1l85, Ln1l85, Sn1l85;
wire Zn1l85, Go1l85, No1l85, Uo1l85, Bp1l85, Ip1l85, Pp1l85, Wp1l85, Dq1l85, Kq1l85;
wire Rq1l85, Yq1l85, Fr1l85, Mr1l85, Tr1l85, As1l85, Hs1l85, Os1l85, Vs1l85, Ct1l85;
wire Jt1l85, Qt1l85, Xt1l85, Eu1l85, Lu1l85, Su1l85, Zu1l85, Gv1l85, Nv1l85, Uv1l85;
wire Bw1l85;
wire [3:0] Iw1l85;
wire [30:2] Nx1l85;
wire [31:0] Sy1l85;
wire [31:0] Tz1l85;
wire [31:0] B12l85;
wire [31:0] J22l85;
wire [8:1] R32l85;
wire [30:0] E52l85;
wire [1:0] M62l85;
wire [23:0] V72l85;
wire [1:0] C92l85;
wire [1:0] Ha2l85;
wire [63:0] Mb2l85;
wire [23:0] Vc2l85;
wire [1:0] Ge2l85;
wire [23:0] Pf2l85;
wire [31:0] Yg2l85;
wire [31:0] Gi2l85;
wire [31:0] Qj2l85;
wire Al2l85, Yl2l85, Wm2l85, Un2l85, So2l85, Qp2l85, Oq2l85, Mr2l85, Ks2l85, It2l85;
wire Gu2l85, Fv2l85, Ew2l85, Dx2l85, Cy2l85, Bz2l85, A03l85, Z03l85, Y13l85, X23l85;
wire W33l85, V43l85, U53l85, T63l85, S73l85, R83l85, Q93l85, Pa3l85, Ob3l85, Nc3l85;
wire Md3l85, Le3l85, Kf3l85, Jg3l85;
reg Ih3l85, Yi3l85, Gk3l85, Vl3l85, Fn3l85, Oo3l85, Yp3l85, Hr3l85, Qs3l85, Fu3l85;
reg Xv3l85, Kx3l85, Vy3l85, I04l85, W14l85, L34l85, Z44l85, O64l85, D84l85, V94l85;
reg Jb4l85, Xc4l85, Pe4l85, Dg4l85, Rh4l85, Fj4l85, Tk4l85, Hm4l85, Zn4l85, Kp4l85;
reg Yq4l85, Os4l85, Du4l85, Sv4l85, Kx4l85, Wy4l85, J05l85, W15l85, K35l85, Z45l85;
reg N65l85, B85l85, Q95l85, Fb5l85, Tc5l85, He5l85, Wf5l85, Lh5l85, Bj5l85, Qk5l85;
reg Fm5l85, Un5l85, Jp5l85, Br5l85, Ps5l85, Du5l85, Ov5l85, Cx5l85, Qy5l85, E06l85;
reg S16l85, K36l85, V46l85, G66l85, V76l85, I96l85, Va6l85, Fc6l85, Vd6l85, Hf6l85;
reg Wg6l85, Li6l85, Ak6l85, Ml6l85, Bn6l85, Po6l85, Dq6l85, Rr6l85, Ft6l85, Tu6l85;
reg Lw6l85, Ux6l85, Jz6l85, Y07l85, N27l85, C47l85, U57l85, F77l85, T87l85, Ja7l85;
reg Yb7l85, Nd7l85, Cf7l85, Rg7l85, Gi7l85, Vj7l85, Kl7l85, Zm7l85, Qo7l85, Hq7l85;
reg Yr7l85, Pt7l85, Gv7l85, Xw7l85, Oy7l85, F08l85, W18l85, N38l85, E58l85, T68l85;
reg I88l85, X98l85, Ib8l85, Xc8l85, Ke8l85, Xf8l85, Kh8l85, Yi8l85, Jk8l85, Xl8l85;
reg Ln8l85, Zo8l85, Nq8l85, Es8l85, Vt8l85, Kv8l85, Zw8l85, Oy8l85, D09l85, V19l85;
reg J39l85, X49l85, L69l85, Z79l85, Q99l85, Eb9l85, Sc9l85, Ge9l85, Uf9l85, Ih9l85;
reg Wi9l85, Kk9l85, Bm9l85, Sn9l85, Ip9l85, Yq9l85, Ns9l85, Cu9l85, Rv9l85, Gx9l85;
reg Xy9l85, O0al85, B2al85, P3al85, F5al85, V6al85, M8al85, Aaal85, Obal85, Cdal85;
reg Qeal85, Hgal85, Yhal85, Mjal85, Alal85, Omal85, Coal85, Qpal85, Eral85, Ssal85;
reg Jual85, Awal85, Pxal85, Ezal85, T0bl85, I2bl85, A4bl85, L5bl85, D7bl85, V8bl85;
reg Kabl85, Zbbl85, Odbl85, Dfbl85, Vgbl85, Kibl85, Zjbl85, Olbl85, Dnbl85, Sobl85;
reg Hqbl85, Wrbl85, Ltbl85, Avbl85, Pwbl85, Eybl85, Tzbl85, I1cl85, A3cl85, P4cl85;
reg E6cl85, T7cl85, I9cl85, Abcl85, Occl85, Cecl85, Qfcl85, Dhcl85, Qicl85, Bkcl85;
reg Nlcl85, Bncl85, Pocl85, Dqcl85, Rrcl85, Gtcl85, Vucl85, Kwcl85, Zxcl85, Nzcl85;
reg Z0dl85, L2dl85, B4dl85, N5dl85, Z6dl85, L8dl85, Cadl85, Ubdl85, Iddl85, Xedl85;
reg Lgdl85, Zhdl85, Njdl85, Bldl85, Pmdl85, Dodl85, Rpdl85, Frdl85, Tsdl85, Hudl85;
reg Wvdl85, Lxdl85, Azdl85, P0el85, E2el85, T3el85, I5el85, W6el85, K8el85, Y9el85;
reg Nbel85, Edel85, Veel85, Mgel85, Diel85, Pjel85, Clel85, Nmel85, Znel85, Kpel85;
reg Vqel85, Gsel85, Rtel85, Cvel85, Nwel85, Yxel85, Kzel85, W0fl85, I2fl85, U3fl85;
reg G5fl85, S6fl85, E8fl85, Q9fl85, Cbfl85, Ocfl85, Aefl85, Mffl85, Ygfl85, Kifl85;
reg Wjfl85, Ilfl85, Wmfl85, Kofl85, Ypfl85, Mrfl85, Atfl85, Oufl85, Cwfl85, Qxfl85;
reg Fzfl85, U0gl85, J2gl85, U3gl85, M5gl85, E7gl85, W8gl85, Kagl85, Ybgl85, Mdgl85;
reg Afgl85, Oggl85, Digl85, Sjgl85, Glgl85, Umgl85, Iogl85, Xpgl85, Mrgl85, Btgl85;
reg Qugl85, Fwgl85, Uxgl85, Izgl85, W0hl85, K2hl85, Y3hl85, N5hl85, C7hl85, R8hl85;
reg Gahl85, Vbhl85, Kdhl85, Zehl85, Nghl85, Bihl85, Qjhl85, Flhl85, Umhl85, Iohl85;
reg Wphl85, Krhl85, Zshl85, Ouhl85, Dwhl85, Sxhl85, Hzhl85, W0il85, K2il85, Y3il85;
reg M5il85, A7il85, P8il85, Eail85, Tbil85, Idil85, Xeil85, Mgil85, Biil85, Pjil85;
reg Dlil85, Smil85, Goil85, Vpil85, Kril85, Zsil85, Ouil85, Dwil85, Sxil85, Hzil85;
reg V0jl85, J2jl85, X3jl85, L5jl85, A7jl85, P8jl85, Eajl85, Tbjl85, Hdjl85, Vejl85;
reg Jgjl85, Yhjl85, Njjl85, Cljl85, Rmjl85, Fojl85, Tpjl85, Hrjl85, Wsjl85, Lujl85;
reg Awjl85, Pxjl85, Ezjl85, S0kl85, G2kl85, U3kl85, I5kl85, X6kl85, M8kl85, Bakl85;
reg Qbkl85, Edkl85, Sekl85, Hgkl85, Whkl85, Kjkl85, Ykkl85, Mmkl85, Bokl85, Qpkl85;
reg Frkl85, Uskl85, Jukl85, Xvkl85, Lxkl85, Zykl85, N0ll85, C2ll85, R3ll85, G5ll85;
reg V6ll85, J8ll85, X9ll85, Mbll85, Bdll85, Pell85, Dgll85, Rhll85, Gjll85, Vkll85;
reg Kmll85, Znll85, Opll85, Drll85, Rsll85, Full85, Tvll85, Hxll85, Wyll85, L0ml85;
reg A2ml85, P3ml85, E5ml85, T6ml85, I8ml85, W9ml85, Kbml85, Zcml85, Oeml85, Dgml85;
reg Rhml85, Fjml85, Tkml85, Imml85, Xnml85, Mpml85, Brml85, Qsml85, Fuml85, Tvml85;
reg Hxml85, Vyml85, J0nl85, Y1nl85, N3nl85, C5nl85, R6nl85, G8nl85, V9nl85, Kbnl85;
reg Ycnl85, Menl85, Bgnl85, Qhnl85, Fjnl85, Tknl85, Hmnl85, Vnnl85, Kpnl85, Zqnl85;
reg Osnl85, Dunl85, Svnl85, Hxnl85, Vynl85, J0ol85, X1ol85, L3ol85, A5ol85, P6ol85;
reg E8ol85, T9ol85, Ibol85, Xcol85, Meol85, Agol85, Ohol85, Djol85, Skol85, Hmol85;
reg Vnol85, Jpol85, Xqol85, Msol85, Buol85, Qvol85, Fxol85, Uyol85, J0pl85, X1pl85;
reg L3pl85, Z4pl85, N6pl85, C8pl85, R9pl85, Gbpl85, Vcpl85, Kepl85, Zfpl85, Ohpl85;
reg Cjpl85, Qkpl85, Fmpl85, Unpl85, Jppl85, Xqpl85, Lspl85, Ztpl85, Ovpl85, Dxpl85;
reg Sypl85, H0ql85, W1ql85, L3ql85, Z4ql85, N6ql85, B8ql85, P9ql85, Ebql85, Tcql85;
reg Ieql85, Xfql85, Mhql85, Bjql85, Qkql85, Emql85, Snql85, Hpql85, Wqql85, Lsql85;
reg Ztql85, Nvql85, Bxql85, Qyql85, F0rl85, U1rl85, J3rl85, Y4rl85, N6rl85, B8rl85;
reg P9rl85, Dbrl85, Rcrl85, Gerl85, Vfrl85, Khrl85, Zirl85, Okrl85, Dmrl85, Snrl85;
reg Gprl85, Uqrl85, Jsrl85, Ytrl85, Nvrl85, Cxrl85, Ryrl85, G0sl85, V1sl85, J3sl85;
reg X4sl85, L6sl85, Z7sl85, N9sl85, Cbsl85, Rcsl85, Gesl85, Vfsl85, Khsl85, Zisl85;
reg Oksl85, Cmsl85, Qnsl85, Epsl85, Sqsl85, Gssl85, Utsl85, Ivsl85, Wwsl85, Kysl85;
reg Yzsl85, M1tl85, A3tl85, O4tl85, C6tl85, Q7tl85, E9tl85, Satl85, Gctl85, Udtl85;
reg Jftl85, Zgtl85, Nitl85, Bktl85, Nltl85, Cntl85, Rotl85, Gqtl85, Vrtl85, Kttl85;
reg Zutl85, Owtl85, Dytl85, Sztl85, H1ul85, W2ul85, L4ul85, A6ul85, P7ul85, F9ul85;
reg Vaul85, Jcul85, Xdul85, Lful85, Zgul85, Piul85, Ekul85, Tlul85, Inul85, Xoul85;
reg Mqul85, Bsul85, Qtul85, Fvul85, Vwul85, Lyul85, B0vl85, R1vl85, H3vl85, X4vl85;
reg N6vl85, D8vl85, T9vl85, Jbvl85, Zcvl85, Pevl85, Fgvl85, Vhvl85, Ljvl85, Blvl85;
reg Rmvl85, Hovl85, Wpvl85, Mrvl85, Atvl85, Ouvl85, Cwvl85, Rxvl85, Izvl85, Y0wl85;
reg O2wl85, F4wl85, W5wl85, N7wl85, E9wl85, Vawl85, Lcwl85, Bewl85, Rfwl85, Hhwl85;
reg Xiwl85, Nkwl85, Dmwl85, Tnwl85, Kpwl85, Brwl85, Sswl85, Juwl85, Awwl85, Rxwl85;
reg Izwl85, Z0xl85, Q2xl85, H4xl85, Y5xl85, P7xl85, G9xl85, Xaxl85, Ocxl85, Fexl85;
reg Wfxl85, Nhxl85, Ejxl85, Vkxl85, Mmxl85, Doxl85, Upxl85, Lrxl85, Dtxl85, Vuxl85;
reg Nwxl85, Fyxl85, Wzxl85, N1yl85, E3yl85, V4yl85, N6yl85, F8yl85, X9yl85, Pbyl85;
reg Gdyl85, Yeyl85, Qgyl85, Iiyl85, Zjyl85, Qlyl85, Hnyl85, Yoyl85, Pqyl85, Gsyl85;
reg Xtyl85, Ovyl85, Fxyl85, Wyyl85, O0zl85, G2zl85, Y3zl85, Q5zl85, I7zl85, A9zl85;
reg Sazl85, Kczl85, Cezl85, Ufzl85, Mhzl85, Ejzl85, Vkzl85, Mmzl85, Dozl85, Upzl85;
reg Lrzl85, Ctzl85, Tuzl85, Kwzl85, Ayzl85, Rzzl85, I10m85, W20m85, K40m85, B60m85;
reg S70m85, I90m85, Ya0m85, Oc0m85, Ee0m85, Pf0m85, Fh0m85, Vi0m85, Lk0m85, Bm0m85;
reg Rn0m85, Hp0m85, Xq0m85, Ns0m85, Du0m85, Tv0m85, Jx0m85, Zy0m85, Q01m85, H21m85;
reg Y31m85, P51m85, G71m85, X81m85, Oa1m85, Fc1m85, Wd1m85, Nf1m85, Eh1m85, Vi1m85;
reg Kk1m85, Zl1m85, On1m85, Dp1m85, Sq1m85, Hs1m85, Wt1m85, Lv1m85, Ax1m85, Py1m85;
reg E02m85, T12m85, I32m85, U42m85, J62m85, Y72m85, M92m85, Ab2m85, Pc2m85, Ee2m85;
reg Tf2m85, Ih2m85, Xi2m85, Mk2m85, Bm2m85, Qn2m85, Fp2m85, Uq2m85, Js2m85, Yt2m85;
reg Nv2m85, Zw2m85, Oy2m85, D03m85, R13m85, F33m85, V43m85, M63m85, D83m85, S93m85;
reg Hb3m85, Wc3m85, Le3m85, Ag3m85, Ph3m85, Ej3m85, Tk3m85, Im3m85, Xn3m85, Mp3m85;
reg Br3m85, Qs3m85, Cu3m85, Rv3m85, Gx3m85, Vy3m85, K04m85, A24m85, R34m85, I54m85;
reg A74m85, S84m85, Ha4m85, Wb4m85, Ld4m85, Af4m85, Pg4m85, Ei4m85, Tj4m85, Il4m85;
reg Xm4m85, Mo4m85, Bq4m85, Qr4m85, Ft4m85, Uu4m85, Jw4m85, Yx4m85, Nz4m85, D15m85;
reg U25m85, L45m85, D65m85, V75m85, K95m85, Za5m85, Oc5m85, De5m85, Sf5m85, Hh5m85;
reg Wi5m85, Lk5m85, Am5m85, Pn5m85, Bp5m85, Qq5m85, Fs5m85, Ut5m85, Jv5m85, Yw5m85;
reg Ny5m85, C06m85, R16m85, G36m85, V46m85, K66m85, Z76m85, O96m85, Db6m85, Sc6m85;
reg He6m85, Wf6m85, Lh6m85, Aj6m85, Pk6m85, Em6m85, Tn6m85, Ip6m85, Xq6m85, Ms6m85;
reg Bu6m85, Qv6m85, Fx6m85, Uy6m85, J07m85, Y17m85, N37m85, E57m85, V67m85, N87m85;
reg Ca7m85, Rb7m85, Gd7m85, Ve7m85, Kg7m85, Zh7m85, Oj7m85, Dl7m85, Sm7m85, Ho7m85;
reg Xp7m85, Mr7m85;
wire [33:0] Dt7m85;
wire [33:0] Tu7m85;

assign hprot_o[1] = 1'b1;
assign hburst_o[2] = 1'b0;
assign hburst_o[1] = 1'b0;
assign hburst_o[0] = 1'b0;
assign hmastlock_o = 1'b0;
assign hsize_o[2] = 1'b0;
assign htrans_o[0] = 1'b0;
assign Ker675 = Ih3l85;
assign vis_tbit_o = Yi3l85;
assign Rpi675 = Gk3l85;
assign C4i675 = Vl3l85;
assign vis_apsr_o[3] = Fn3l85;
assign Gvo675 = Oo3l85;
assign vis_apsr_o[1] = Yp3l85;
assign vis_apsr_o[2] = Hr3l85;
assign Krm675 = Qs3l85;
assign Gi2l85[30] = Fu3l85;
assign Hph675 = Xv3l85;
assign Bvh675 = Kx3l85;
assign O4p675 = Vy3l85;
assign Iw1l85[3] = I04l85;
assign vis_r7_o[23] = W14l85;
assign C92l85[1] = L34l85;
assign vis_r7_o[31] = Z44l85;
assign vis_r0_o[31] = O64l85;
assign Gi2l85[31] = D84l85;
assign vis_r7_o[7] = V94l85;
assign vis_r0_o[7] = Jb4l85;
assign Gi2l85[15] = Xc4l85;
assign Z9n675 = Pe4l85;
assign T7i675 = Dg4l85;
assign Hsi675 = Rh4l85;
assign vis_r7_o[1] = Fj4l85;
assign vis_r0_o[1] = Tk4l85;
assign Gi2l85[25] = Hm4l85;
assign vis_ipsr_o[1] = Zn4l85;
assign Mml675 = Kp4l85;
assign M62l85[1] = Yq4l85;
assign vis_r7_o[14] = Os4l85;
assign vis_psp_o[12] = Du4l85;
assign Gi2l85[14] = Sv4l85;
assign vis_pc_o[29] = Kx4l85;
assign Vxo675 = Wy4l85;
assign Ezo675 = J05l85;
assign Iw1l85[0] = W15l85;
assign vis_r5_o[31] = K35l85;
assign vis_r5_o[7] = Z45l85;
assign vis_r5_o[1] = N65l85;
assign vis_r5_o[14] = B85l85;
assign vis_r1_o[31] = Q95l85;
assign vis_r1_o[7] = Fb5l85;
assign vis_r1_o[1] = Tc5l85;
assign vis_r1_o[14] = He5l85;
assign vis_r1_o[23] = Wf5l85;
assign O8r675 = Lh5l85;
assign vis_r1_o[24] = Bj5l85;
assign vis_r5_o[24] = Qk5l85;
assign vis_r7_o[24] = Fm5l85;
assign vis_psp_o[22] = Un5l85;
assign Gi2l85[24] = Jp5l85;
assign Tcn675 = Br5l85;
assign Pui675 = Ps5l85;
assign vis_control_o = Du5l85;
assign vis_r1_o[2] = Ov5l85;
assign vis_r5_o[2] = Cx5l85;
assign vis_r7_o[2] = Qy5l85;
assign vis_psp_o[0] = E06l85;
assign Gi2l85[10] = S16l85;
assign vis_ipsr_o[2] = K36l85;
assign vis_pc_o[0] = V46l85;
assign Gwh675 = G66l85;
assign F3p675 = V76l85;
assign W1p675 = I96l85;
assign X5p675 = Va6l85;
assign J7p675 = Fc6l85;
assign Cep675 = Vd6l85;
assign Jwn675 = Hf6l85;
assign Ntn675 = Wg6l85;
assign Yun675 = Li6l85;
assign Nvm675 = Ak6l85;
assign Zqi675 = Ml6l85;
assign Xwi675 = Bn6l85;
assign vis_r1_o[4] = Po6l85;
assign vis_r5_o[4] = Dq6l85;
assign vis_r7_o[4] = Rr6l85;
assign vis_psp_o[2] = Ft6l85;
assign Gi2l85[20] = Tu6l85;
assign vis_apsr_o[0] = Lw6l85;
assign vis_r5_o[28] = Ux6l85;
assign vis_r7_o[28] = Jz6l85;
assign vis_r1_o[28] = Y07l85;
assign vis_r0_o[28] = N27l85;
assign Gi2l85[28] = C47l85;
assign vis_ipsr_o[4] = U57l85;
assign Qql675 = F77l85;
assign Aar675 = T87l85;
assign vis_r1_o[15] = Ja7l85;
assign vis_r5_o[15] = Yb7l85;
assign vis_r7_o[15] = Nd7l85;
assign vis_r1_o[30] = Cf7l85;
assign vis_r5_o[30] = Rg7l85;
assign vis_r7_o[30] = Gi7l85;
assign vis_psp_o[28] = Vj7l85;
assign Lnh675 = Kl7l85;
assign Mb2l85[58] = Zm7l85;
assign Mb2l85[59] = Qo7l85;
assign Mb2l85[61] = Hq7l85;
assign Mb2l85[62] = Yr7l85;
assign Mb2l85[63] = Pt7l85;
assign Mb2l85[26] = Gv7l85;
assign Mb2l85[27] = Xw7l85;
assign Mb2l85[29] = Oy7l85;
assign Mb2l85[30] = F08l85;
assign Mb2l85[31] = W18l85;
assign Gi2l85[9] = N38l85;
assign vis_r1_o[25] = E58l85;
assign vis_r5_o[25] = T68l85;
assign vis_r7_o[25] = I88l85;
assign vis_ipsr_o[3] = X98l85;
assign Jqh675 = Ib8l85;
assign Rto675 = Xc8l85;
assign N0p675 = Ke8l85;
assign Mwo675 = Xf8l85;
assign E0i675 = Kh8l85;
assign vis_primask_o = Yi8l85;
assign vis_r5_o[0] = Jk8l85;
assign vis_r7_o[0] = Xl8l85;
assign vis_r1_o[0] = Ln8l85;
assign vis_r0_o[0] = Zo8l85;
assign Qj2l85[0] = Nq8l85;
assign Gi2l85[0] = Es8l85;
assign vis_r1_o[16] = Vt8l85;
assign vis_r5_o[16] = Kv8l85;
assign vis_r7_o[16] = Zw8l85;
assign vis_psp_o[14] = Oy8l85;
assign Gi2l85[16] = D09l85;
assign vis_r1_o[8] = V19l85;
assign vis_r5_o[8] = J39l85;
assign vis_r7_o[8] = X49l85;
assign vis_psp_o[6] = L69l85;
assign Gi2l85[8] = Z79l85;
assign Jbn675 = Q99l85;
assign A9i675 = Eb9l85;
assign Lti675 = Sc9l85;
assign vis_r1_o[3] = Ge9l85;
assign vis_r5_o[3] = Uf9l85;
assign vis_r7_o[3] = Ih9l85;
assign vis_psp_o[1] = Wi9l85;
assign Pf2l85[19] = Kk9l85;
assign V72l85[19] = Bm9l85;
assign V72l85[0] = Sn9l85;
assign V72l85[1] = Ip9l85;
assign vis_r1_o[17] = Yq9l85;
assign vis_r5_o[17] = Ns9l85;
assign vis_r7_o[17] = Cu9l85;
assign vis_psp_o[15] = Rv9l85;
assign Pf2l85[17] = Gx9l85;
assign V72l85[17] = Xy9l85;
assign N6i675 = O0al85;
assign Oxl675 = B2al85;
assign Pf2l85[9] = P3al85;
assign V72l85[9] = F5al85;
assign V72l85[22] = V6al85;
assign vis_r1_o[6] = M8al85;
assign vis_r5_o[6] = Aaal85;
assign vis_r7_o[6] = Obal85;
assign vis_psp_o[4] = Cdal85;
assign Mb2l85[60] = Qeal85;
assign Mb2l85[28] = Hgal85;
assign C92l85[0] = Yhal85;
assign Xgn675 = Mjal85;
assign Byi675 = Alal85;
assign vis_r1_o[5] = Omal85;
assign vis_r5_o[5] = Coal85;
assign vis_r7_o[5] = Qpal85;
assign vis_psp_o[3] = Eral85;
assign Pf2l85[21] = Ssal85;
assign V72l85[21] = Jual85;
assign vis_r1_o[29] = Awal85;
assign vis_r5_o[29] = Pxal85;
assign vis_r7_o[29] = Ezal85;
assign vis_psp_o[27] = T0bl85;
assign Gi2l85[29] = I2bl85;
assign vis_ipsr_o[5] = A4bl85;
assign Qj2l85[11] = L5bl85;
assign Gi2l85[11] = D7bl85;
assign vis_r1_o[27] = V8bl85;
assign vis_r5_o[27] = Kabl85;
assign vis_r7_o[27] = Zbbl85;
assign vis_psp_o[25] = Odbl85;
assign Gi2l85[27] = Dfbl85;
assign vis_r1_o[19] = Vgbl85;
assign vis_r5_o[19] = Kibl85;
assign vis_r7_o[19] = Zjbl85;
assign vis_r1_o[20] = Olbl85;
assign vis_r5_o[20] = Dnbl85;
assign vis_r7_o[20] = Sobl85;
assign vis_r1_o[21] = Hqbl85;
assign vis_r5_o[21] = Wrbl85;
assign vis_r7_o[21] = Ltbl85;
assign vis_r1_o[26] = Avbl85;
assign vis_r5_o[26] = Pwbl85;
assign vis_r7_o[26] = Eybl85;
assign vis_psp_o[24] = Tzbl85;
assign Gi2l85[26] = I1cl85;
assign vis_r1_o[18] = A3cl85;
assign vis_r5_o[18] = P4cl85;
assign vis_r7_o[18] = E6cl85;
assign vis_psp_o[16] = T7cl85;
assign Gi2l85[18] = I9cl85;
assign Nfn675 = Abcl85;
assign Den675 = Occl85;
assign P8n675 = Cecl85;
assign Iso675 = Qfcl85;
assign Lrh675 = Dhcl85;
assign vis_ipsr_o[0] = Qicl85;
assign Ogp675 = Bkcl85;
assign Hin675 = Nlcl85;
assign Rjn675 = Bncl85;
assign Bln675 = Pocl85;
assign Lmn675 = Dqcl85;
assign Vnn675 = Rrcl85;
assign Gpn675 = Gtcl85;
assign Rqn675 = Vucl85;
assign Csn675 = Kwcl85;
assign Tvi675 = Zxcl85;
assign vis_pc_o[21] = Nzcl85;
assign vis_pc_o[30] = Z0dl85;
assign Ycr675 = L2dl85;
assign Skp675 = B4dl85;
assign Wcp675 = N5dl85;
assign Ifp675 = Z6dl85;
assign Doh675 = L8dl85;
assign N1j675 = Cadl85;
assign Plo675 = Ubdl85;
assign Eko675 = Iddl85;
assign Uxn675 = Xedl85;
assign Ezn675 = Lgdl85;
assign O0o675 = Zhdl85;
assign Y1o675 = Njdl85;
assign I3o675 = Bldl85;
assign S4o675 = Pmdl85;
assign C6o675 = Dodl85;
assign M7o675 = Rpdl85;
assign W8o675 = Frdl85;
assign Gao675 = Tsdl85;
assign Qbo675 = Hudl85;
assign Bdo675 = Wvdl85;
assign Meo675 = Lxdl85;
assign Xfo675 = Azdl85;
assign Iho675 = P0el85;
assign Tio675 = E2el85;
assign Joi675 = T3el85;
assign Iw1l85[1] = I5el85;
assign V8p675 = W6el85;
assign Oxh675 = K8el85;
assign Nbp675 = Y9el85;
assign Mb2l85[56] = Nbel85;
assign Mb2l85[24] = Edel85;
assign Mb2l85[57] = Veel85;
assign Mb2l85[25] = Mgel85;
assign Tth675 = Diel85;
assign G5i675 = Pjel85;
assign vis_pc_o[1] = Clel85;
assign Lsh675 = Nmel85;
assign vis_pc_o[2] = Znel85;
assign vis_pc_o[3] = Kpel85;
assign vis_pc_o[4] = Vqel85;
assign vis_pc_o[5] = Gsel85;
assign vis_pc_o[6] = Rtel85;
assign vis_pc_o[7] = Cvel85;
assign vis_pc_o[8] = Nwel85;
assign vis_pc_o[13] = Yxel85;
assign vis_pc_o[14] = Kzel85;
assign vis_pc_o[15] = W0fl85;
assign vis_pc_o[16] = I2fl85;
assign vis_pc_o[17] = U3fl85;
assign vis_pc_o[18] = G5fl85;
assign vis_pc_o[19] = S6fl85;
assign vis_pc_o[20] = E8fl85;
assign vis_pc_o[23] = Q9fl85;
assign vis_pc_o[24] = Cbfl85;
assign vis_pc_o[25] = Ocfl85;
assign vis_pc_o[26] = Aefl85;
assign vis_pc_o[27] = Mffl85;
assign vis_pc_o[28] = Ygfl85;
assign Spo675 = Kifl85;
assign Aro675 = Wjfl85;
assign Hai675 = Ilfl85;
assign Obi675 = Wmfl85;
assign Vci675 = Kofl85;
assign Cei675 = Ypfl85;
assign Jfi675 = Mrfl85;
assign Qgi675 = Atfl85;
assign Xhi675 = Oufl85;
assign Eji675 = Cwfl85;
assign Lki675 = Qxfl85;
assign Tli675 = Fzfl85;
assign Bni675 = U0gl85;
assign Gum675 = J2gl85;
assign R2j675 = U3gl85;
assign V3j675 = M5gl85;
assign A5j675 = E7gl85;
assign M1i675 = W8gl85;
assign Fzi675 = Kagl85;
assign J0j675 = Ybgl85;
assign U2i675 = Mdgl85;
assign Iw1l85[2] = Afgl85;
assign vis_r6_o[31] = Oggl85;
assign vis_r6_o[28] = Digl85;
assign vis_r6_o[7] = Sjgl85;
assign vis_r6_o[1] = Glgl85;
assign vis_r6_o[0] = Umgl85;
assign vis_r6_o[30] = Iogl85;
assign vis_r6_o[29] = Xpgl85;
assign vis_r6_o[27] = Mrgl85;
assign vis_r6_o[26] = Btgl85;
assign vis_r6_o[25] = Qugl85;
assign vis_r6_o[24] = Fwgl85;
assign vis_r6_o[6] = Uxgl85;
assign vis_r6_o[5] = Izgl85;
assign vis_r6_o[4] = W0hl85;
assign vis_r6_o[3] = K2hl85;
assign vis_r6_o[21] = Y3hl85;
assign vis_r6_o[20] = N5hl85;
assign vis_r6_o[19] = C7hl85;
assign vis_r6_o[18] = R8hl85;
assign vis_r6_o[17] = Gahl85;
assign vis_r6_o[16] = Vbhl85;
assign vis_r6_o[14] = Kdhl85;
assign vis_r6_o[2] = Zehl85;
assign vis_r6_o[8] = Nghl85;
assign vis_r6_o[15] = Bihl85;
assign vis_r4_o[31] = Qjhl85;
assign vis_r4_o[28] = Flhl85;
assign vis_r4_o[7] = Umhl85;
assign vis_r4_o[1] = Iohl85;
assign vis_r4_o[0] = Wphl85;
assign vis_r4_o[30] = Krhl85;
assign vis_r4_o[29] = Zshl85;
assign vis_r4_o[27] = Ouhl85;
assign vis_r4_o[26] = Dwhl85;
assign vis_r4_o[25] = Sxhl85;
assign vis_r4_o[24] = Hzhl85;
assign vis_r4_o[6] = W0il85;
assign vis_r4_o[5] = K2il85;
assign vis_r4_o[4] = Y3il85;
assign vis_r4_o[3] = M5il85;
assign vis_r4_o[21] = A7il85;
assign vis_r4_o[20] = P8il85;
assign vis_r4_o[19] = Eail85;
assign vis_r4_o[18] = Tbil85;
assign vis_r4_o[17] = Idil85;
assign vis_r4_o[16] = Xeil85;
assign vis_r4_o[14] = Mgil85;
assign vis_r4_o[2] = Biil85;
assign vis_r4_o[8] = Pjil85;
assign vis_r4_o[15] = Dlil85;
assign vis_msp_o[5] = Smil85;
assign vis_msp_o[26] = Goil85;
assign vis_msp_o[29] = Vpil85;
assign vis_msp_o[28] = Kril85;
assign vis_msp_o[27] = Zsil85;
assign vis_msp_o[25] = Ouil85;
assign vis_msp_o[24] = Dwil85;
assign vis_msp_o[22] = Sxil85;
assign vis_msp_o[4] = Hzil85;
assign vis_msp_o[3] = V0jl85;
assign vis_msp_o[2] = J2jl85;
assign vis_msp_o[1] = X3jl85;
assign vis_msp_o[16] = L5jl85;
assign vis_msp_o[15] = A7jl85;
assign vis_msp_o[14] = P8jl85;
assign vis_msp_o[12] = Eajl85;
assign vis_msp_o[0] = Tbjl85;
assign vis_msp_o[6] = Hdjl85;
assign vis_psp_o[5] = Vejl85;
assign vis_psp_o[26] = Jgjl85;
assign vis_psp_o[29] = Yhjl85;
assign vis_r12_o[31] = Njjl85;
assign vis_r12_o[28] = Cljl85;
assign vis_r12_o[7] = Rmjl85;
assign vis_r12_o[1] = Fojl85;
assign vis_r12_o[0] = Tpjl85;
assign vis_r12_o[30] = Hrjl85;
assign vis_r12_o[29] = Wsjl85;
assign vis_r12_o[27] = Lujl85;
assign vis_r12_o[26] = Awjl85;
assign vis_r12_o[24] = Pxjl85;
assign vis_r12_o[6] = Ezjl85;
assign vis_r12_o[5] = S0kl85;
assign vis_r12_o[4] = G2kl85;
assign vis_r12_o[3] = U3kl85;
assign vis_r12_o[18] = I5kl85;
assign vis_r12_o[17] = X6kl85;
assign vis_r12_o[16] = M8kl85;
assign vis_r12_o[14] = Bakl85;
assign vis_r12_o[2] = Qbkl85;
assign vis_r12_o[8] = Edkl85;
assign vis_r14_o[31] = Sekl85;
assign vis_r14_o[28] = Hgkl85;
assign vis_r14_o[7] = Whkl85;
assign vis_r14_o[1] = Kjkl85;
assign vis_r14_o[0] = Ykkl85;
assign vis_r14_o[30] = Mmkl85;
assign vis_r14_o[29] = Bokl85;
assign vis_r14_o[27] = Qpkl85;
assign vis_r14_o[26] = Frkl85;
assign vis_r14_o[24] = Uskl85;
assign vis_r14_o[6] = Jukl85;
assign vis_r14_o[5] = Xvkl85;
assign vis_r14_o[4] = Lxkl85;
assign vis_r14_o[3] = Zykl85;
assign vis_r14_o[18] = N0ll85;
assign vis_r14_o[17] = C2ll85;
assign vis_r14_o[16] = R3ll85;
assign vis_r14_o[14] = G5ll85;
assign vis_r14_o[2] = V6ll85;
assign vis_r14_o[8] = J8ll85;
assign vis_r11_o[31] = X9ll85;
assign vis_r11_o[28] = Mbll85;
assign vis_r11_o[7] = Bdll85;
assign vis_r11_o[1] = Pell85;
assign vis_r11_o[0] = Dgll85;
assign vis_r11_o[30] = Rhll85;
assign vis_r11_o[29] = Gjll85;
assign vis_r11_o[27] = Vkll85;
assign vis_r11_o[26] = Kmll85;
assign vis_r11_o[25] = Znll85;
assign vis_r11_o[24] = Opll85;
assign vis_r11_o[6] = Drll85;
assign vis_r11_o[5] = Rsll85;
assign vis_r11_o[4] = Full85;
assign vis_r11_o[3] = Tvll85;
assign vis_r11_o[21] = Hxll85;
assign vis_r11_o[20] = Wyll85;
assign vis_r11_o[19] = L0ml85;
assign vis_r11_o[18] = A2ml85;
assign vis_r11_o[17] = P3ml85;
assign vis_r11_o[16] = E5ml85;
assign vis_r11_o[14] = T6ml85;
assign vis_r11_o[2] = I8ml85;
assign vis_r11_o[8] = W9ml85;
assign vis_r11_o[15] = Kbml85;
assign vis_r10_o[31] = Zcml85;
assign vis_r10_o[28] = Oeml85;
assign vis_r10_o[7] = Dgml85;
assign vis_r10_o[1] = Rhml85;
assign vis_r10_o[0] = Fjml85;
assign vis_r10_o[30] = Tkml85;
assign vis_r10_o[29] = Imml85;
assign vis_r10_o[27] = Xnml85;
assign vis_r10_o[26] = Mpml85;
assign vis_r10_o[25] = Brml85;
assign vis_r10_o[24] = Qsml85;
assign vis_r10_o[6] = Fuml85;
assign vis_r10_o[5] = Tvml85;
assign vis_r10_o[4] = Hxml85;
assign vis_r10_o[3] = Vyml85;
assign vis_r10_o[21] = J0nl85;
assign vis_r10_o[20] = Y1nl85;
assign vis_r10_o[19] = N3nl85;
assign vis_r10_o[18] = C5nl85;
assign vis_r10_o[17] = R6nl85;
assign vis_r10_o[16] = G8nl85;
assign vis_r10_o[14] = V9nl85;
assign vis_r10_o[2] = Kbnl85;
assign vis_r10_o[8] = Ycnl85;
assign vis_r10_o[15] = Menl85;
assign vis_r9_o[31] = Bgnl85;
assign vis_r9_o[28] = Qhnl85;
assign vis_r9_o[7] = Fjnl85;
assign vis_r9_o[1] = Tknl85;
assign vis_r9_o[0] = Hmnl85;
assign vis_r9_o[30] = Vnnl85;
assign vis_r9_o[29] = Kpnl85;
assign vis_r9_o[27] = Zqnl85;
assign vis_r9_o[26] = Osnl85;
assign vis_r9_o[25] = Dunl85;
assign vis_r9_o[24] = Svnl85;
assign vis_r9_o[6] = Hxnl85;
assign vis_r9_o[5] = Vynl85;
assign vis_r9_o[4] = J0ol85;
assign vis_r9_o[3] = X1ol85;
assign vis_r9_o[21] = L3ol85;
assign vis_r9_o[20] = A5ol85;
assign vis_r9_o[19] = P6ol85;
assign vis_r9_o[18] = E8ol85;
assign vis_r9_o[17] = T9ol85;
assign vis_r9_o[16] = Ibol85;
assign vis_r9_o[14] = Xcol85;
assign vis_r9_o[2] = Meol85;
assign vis_r9_o[8] = Agol85;
assign vis_r9_o[15] = Ohol85;
assign vis_r8_o[31] = Djol85;
assign vis_r8_o[28] = Skol85;
assign vis_r8_o[7] = Hmol85;
assign vis_r8_o[1] = Vnol85;
assign vis_r8_o[0] = Jpol85;
assign vis_r8_o[30] = Xqol85;
assign vis_r8_o[29] = Msol85;
assign vis_r8_o[27] = Buol85;
assign vis_r8_o[26] = Qvol85;
assign vis_r8_o[25] = Fxol85;
assign vis_r8_o[24] = Uyol85;
assign vis_r8_o[6] = J0pl85;
assign vis_r8_o[5] = X1pl85;
assign vis_r8_o[4] = L3pl85;
assign vis_r8_o[3] = Z4pl85;
assign vis_r8_o[21] = N6pl85;
assign vis_r8_o[20] = C8pl85;
assign vis_r8_o[19] = R9pl85;
assign vis_r8_o[18] = Gbpl85;
assign vis_r8_o[17] = Vcpl85;
assign vis_r8_o[16] = Kepl85;
assign vis_r8_o[14] = Zfpl85;
assign vis_r8_o[2] = Ohpl85;
assign vis_r8_o[8] = Cjpl85;
assign vis_r8_o[15] = Qkpl85;
assign vis_r3_o[31] = Fmpl85;
assign vis_r3_o[28] = Unpl85;
assign vis_r3_o[7] = Jppl85;
assign vis_r3_o[1] = Xqpl85;
assign vis_r3_o[0] = Lspl85;
assign vis_r3_o[30] = Ztpl85;
assign vis_r3_o[29] = Ovpl85;
assign vis_r3_o[27] = Dxpl85;
assign vis_r3_o[26] = Sypl85;
assign vis_r3_o[25] = H0ql85;
assign vis_r3_o[24] = W1ql85;
assign vis_r3_o[6] = L3ql85;
assign vis_r3_o[5] = Z4ql85;
assign vis_r3_o[4] = N6ql85;
assign vis_r3_o[3] = B8ql85;
assign vis_r3_o[21] = P9ql85;
assign vis_r3_o[20] = Ebql85;
assign vis_r3_o[19] = Tcql85;
assign vis_r3_o[18] = Ieql85;
assign vis_r3_o[17] = Xfql85;
assign vis_r3_o[16] = Mhql85;
assign vis_r3_o[14] = Bjql85;
assign vis_r3_o[2] = Qkql85;
assign vis_r3_o[8] = Emql85;
assign vis_r3_o[15] = Snql85;
assign vis_r2_o[31] = Hpql85;
assign vis_r2_o[28] = Wqql85;
assign vis_r2_o[7] = Lsql85;
assign vis_r2_o[1] = Ztql85;
assign vis_r2_o[0] = Nvql85;
assign vis_r2_o[30] = Bxql85;
assign vis_r2_o[29] = Qyql85;
assign vis_r2_o[27] = F0rl85;
assign vis_r2_o[26] = U1rl85;
assign vis_r2_o[25] = J3rl85;
assign vis_r2_o[24] = Y4rl85;
assign vis_r2_o[6] = N6rl85;
assign vis_r2_o[5] = B8rl85;
assign vis_r2_o[4] = P9rl85;
assign vis_r2_o[3] = Dbrl85;
assign vis_r2_o[21] = Rcrl85;
assign vis_r2_o[20] = Gerl85;
assign vis_r2_o[19] = Vfrl85;
assign vis_r2_o[18] = Khrl85;
assign vis_r2_o[17] = Zirl85;
assign vis_r2_o[16] = Okrl85;
assign vis_r2_o[14] = Dmrl85;
assign vis_r2_o[2] = Snrl85;
assign vis_r2_o[8] = Gprl85;
assign vis_r2_o[15] = Uqrl85;
assign vis_r0_o[30] = Jsrl85;
assign vis_r0_o[29] = Ytrl85;
assign vis_r0_o[27] = Nvrl85;
assign vis_r0_o[26] = Cxrl85;
assign vis_r0_o[25] = Ryrl85;
assign vis_r0_o[24] = G0sl85;
assign vis_r0_o[6] = V1sl85;
assign vis_r0_o[5] = J3sl85;
assign vis_r0_o[4] = X4sl85;
assign vis_r0_o[3] = L6sl85;
assign Gpl675 = Z7sl85;
assign vis_r0_o[21] = N9sl85;
assign vis_r0_o[20] = Cbsl85;
assign vis_r0_o[19] = Rcsl85;
assign vis_r0_o[18] = Gesl85;
assign vis_r0_o[17] = Vfsl85;
assign vis_r0_o[16] = Khsl85;
assign vis_r0_o[14] = Zisl85;
assign vis_r0_o[2] = Oksl85;
assign Wnl675 = Cmsl85;
assign vis_r0_o[9] = Qnsl85;
assign vis_r1_o[9] = Epsl85;
assign vis_r2_o[9] = Sqsl85;
assign vis_r3_o[9] = Gssl85;
assign vis_r8_o[9] = Utsl85;
assign vis_r9_o[9] = Ivsl85;
assign vis_r10_o[9] = Wwsl85;
assign vis_r11_o[9] = Kysl85;
assign vis_r4_o[9] = Yzsl85;
assign vis_r5_o[9] = M1tl85;
assign vis_r6_o[9] = A3tl85;
assign vis_r7_o[9] = O4tl85;
assign vis_r12_o[9] = C6tl85;
assign vis_r14_o[9] = Q7tl85;
assign vis_msp_o[7] = E9tl85;
assign vis_psp_o[7] = Satl85;
assign vis_r0_o[8] = Gctl85;
assign vis_r0_o[15] = Udtl85;
assign M62l85[0] = Jftl85;
assign Cll675 = Zgtl85;
assign Wyh675 = Nitl85;
assign vis_pc_o[22] = Bktl85;
assign vis_r0_o[23] = Nltl85;
assign vis_r2_o[23] = Cntl85;
assign vis_r3_o[23] = Rotl85;
assign vis_r8_o[23] = Gqtl85;
assign vis_r9_o[23] = Vrtl85;
assign vis_r10_o[23] = Kttl85;
assign vis_r11_o[23] = Zutl85;
assign vis_r4_o[23] = Owtl85;
assign vis_r5_o[23] = Dytl85;
assign vis_r6_o[23] = Sztl85;
assign vis_r12_o[23] = H1ul85;
assign vis_r14_o[23] = W2ul85;
assign vis_msp_o[21] = L4ul85;
assign vis_psp_o[21] = A6ul85;
assign Ge2l85[0] = P7ul85;
assign Ge2l85[1] = F9ul85;
assign Asl675 = Vaul85;
assign Ktl675 = Jcul85;
assign Uul675 = Xdul85;
assign Ewl675 = Lful85;
assign Mbr675 = Zgul85;
assign Yg2l85[1] = Piul85;
assign Yg2l85[3] = Ekul85;
assign Yg2l85[4] = Tlul85;
assign Yg2l85[5] = Inul85;
assign Yg2l85[6] = Xoul85;
assign Yg2l85[7] = Mqul85;
assign Yg2l85[8] = Bsul85;
assign Yg2l85[9] = Qtul85;
assign Yg2l85[10] = Fvul85;
assign Yg2l85[14] = Vwul85;
assign Yg2l85[15] = Lyul85;
assign Yg2l85[16] = B0vl85;
assign Yg2l85[17] = R1vl85;
assign Yg2l85[18] = H3vl85;
assign Yg2l85[19] = X4vl85;
assign Yg2l85[20] = N6vl85;
assign Yg2l85[21] = D8vl85;
assign Yg2l85[22] = T9vl85;
assign Yg2l85[23] = Jbvl85;
assign Yg2l85[24] = Zcvl85;
assign Yg2l85[25] = Pevl85;
assign Yg2l85[26] = Fgvl85;
assign Yg2l85[27] = Vhvl85;
assign Yg2l85[28] = Ljvl85;
assign Yg2l85[29] = Blvl85;
assign Yg2l85[30] = Rmvl85;
assign Yg2l85[0] = Hovl85;
assign Yg2l85[31] = Wpvl85;
assign Ha2l85[0] = Mrvl85;
assign Ha2l85[1] = Atvl85;
assign Fap675 = Ouvl85;
assign Yg2l85[2] = Cwvl85;
assign Mb2l85[12] = Rxvl85;
assign Mb2l85[8] = Izvl85;
assign Mb2l85[9] = Y0wl85;
assign Mb2l85[10] = O2wl85;
assign Mb2l85[11] = F4wl85;
assign Mb2l85[13] = W5wl85;
assign Mb2l85[14] = N7wl85;
assign Mb2l85[15] = E9wl85;
assign Mb2l85[4] = Vawl85;
assign Mb2l85[0] = Lcwl85;
assign Mb2l85[1] = Bewl85;
assign Mb2l85[2] = Rfwl85;
assign Mb2l85[3] = Hhwl85;
assign Mb2l85[5] = Xiwl85;
assign Mb2l85[6] = Nkwl85;
assign Mb2l85[7] = Dmwl85;
assign Mb2l85[44] = Tnwl85;
assign Mb2l85[40] = Kpwl85;
assign Mb2l85[41] = Brwl85;
assign Mb2l85[42] = Sswl85;
assign Mb2l85[43] = Juwl85;
assign Mb2l85[45] = Awwl85;
assign Mb2l85[46] = Rxwl85;
assign Mb2l85[47] = Izwl85;
assign Mb2l85[36] = Z0xl85;
assign Mb2l85[32] = Q2xl85;
assign Mb2l85[33] = H4xl85;
assign Mb2l85[34] = Y5xl85;
assign Mb2l85[35] = P7xl85;
assign Mb2l85[37] = G9xl85;
assign Mb2l85[38] = Xaxl85;
assign Mb2l85[39] = Ocxl85;
assign Mb2l85[20] = Fexl85;
assign Mb2l85[16] = Wfxl85;
assign Mb2l85[17] = Nhxl85;
assign Mb2l85[18] = Ejxl85;
assign Mb2l85[19] = Vkxl85;
assign Mb2l85[21] = Mmxl85;
assign Mb2l85[22] = Doxl85;
assign Mb2l85[23] = Upxl85;
assign Qj2l85[30] = Lrxl85;
assign Qj2l85[16] = Dtxl85;
assign Qj2l85[17] = Vuxl85;
assign Gi2l85[17] = Nwxl85;
assign Qj2l85[1] = Fyxl85;
assign Gi2l85[1] = Wzxl85;
assign Qj2l85[2] = N1yl85;
assign Gi2l85[2] = E3yl85;
assign Qj2l85[24] = V4yl85;
assign Qj2l85[26] = N6yl85;
assign Qj2l85[27] = F8yl85;
assign Qj2l85[28] = X9yl85;
assign Qj2l85[8] = Pbyl85;
assign Qj2l85[10] = Gdyl85;
assign Qj2l85[14] = Yeyl85;
assign Qj2l85[15] = Qgyl85;
assign Qj2l85[3] = Iiyl85;
assign Gi2l85[3] = Zjyl85;
assign Qj2l85[4] = Qlyl85;
assign Gi2l85[4] = Hnyl85;
assign Qj2l85[5] = Yoyl85;
assign Gi2l85[5] = Pqyl85;
assign Qj2l85[6] = Gsyl85;
assign Gi2l85[6] = Xtyl85;
assign Qj2l85[7] = Ovyl85;
assign Gi2l85[7] = Fxyl85;
assign Qj2l85[20] = Wyyl85;
assign Qj2l85[21] = O0zl85;
assign Gi2l85[21] = G2zl85;
assign Qj2l85[22] = Y3zl85;
assign Gi2l85[22] = Q5zl85;
assign Qj2l85[23] = I7zl85;
assign Gi2l85[23] = A9zl85;
assign Qj2l85[18] = Sazl85;
assign Qj2l85[19] = Kczl85;
assign Gi2l85[19] = Cezl85;
assign Qj2l85[29] = Ufzl85;
assign Qj2l85[31] = Mhzl85;
assign Mb2l85[52] = Ejzl85;
assign Mb2l85[48] = Vkzl85;
assign Mb2l85[49] = Mmzl85;
assign Mb2l85[50] = Dozl85;
assign Mb2l85[51] = Upzl85;
assign Mb2l85[53] = Lrzl85;
assign Mb2l85[54] = Ctzl85;
assign Mb2l85[55] = Tuzl85;
assign S5r675 = Kwzl85;
assign F4r675 = Ayzl85;
assign S2r675 = Rzzl85;
assign E7r675 = I10m85;
assign I1r675 = W20m85;
assign Pf2l85[22] = K40m85;
assign Pf2l85[23] = B60m85;
assign Pf2l85[0] = S70m85;
assign Pf2l85[1] = I90m85;
assign Pf2l85[2] = Ya0m85;
assign V72l85[2] = Oc0m85;
assign vis_pc_o[9] = Ee0m85;
assign Pf2l85[3] = Pf0m85;
assign V72l85[3] = Fh0m85;
assign Pf2l85[4] = Vi0m85;
assign V72l85[4] = Lk0m85;
assign Pf2l85[5] = Bm0m85;
assign V72l85[5] = Rn0m85;
assign Pf2l85[6] = Hp0m85;
assign V72l85[6] = Xq0m85;
assign Pf2l85[7] = Ns0m85;
assign V72l85[7] = Du0m85;
assign Pf2l85[8] = Tv0m85;
assign V72l85[8] = Jx0m85;
assign Pf2l85[10] = Zy0m85;
assign V72l85[10] = Q01m85;
assign Pf2l85[14] = H21m85;
assign V72l85[14] = Y31m85;
assign Pf2l85[15] = P51m85;
assign V72l85[15] = G71m85;
assign Pf2l85[16] = X81m85;
assign V72l85[16] = Oa1m85;
assign Pf2l85[18] = Fc1m85;
assign V72l85[18] = Wd1m85;
assign Pf2l85[20] = Nf1m85;
assign V72l85[20] = Eh1m85;
assign Yyl675 = Vi1m85;
assign vis_r0_o[10] = Kk1m85;
assign vis_r1_o[10] = Zl1m85;
assign vis_r2_o[10] = On1m85;
assign vis_r3_o[10] = Dp1m85;
assign vis_r8_o[10] = Sq1m85;
assign vis_r9_o[10] = Hs1m85;
assign vis_r10_o[10] = Wt1m85;
assign vis_r11_o[10] = Lv1m85;
assign vis_r4_o[10] = Ax1m85;
assign vis_r5_o[10] = Py1m85;
assign vis_r6_o[10] = E02m85;
assign vis_r7_o[10] = T12m85;
assign vis_pc_o[10] = I32m85;
assign vis_r12_o[10] = U42m85;
assign vis_r14_o[10] = J62m85;
assign vis_msp_o[8] = Y72m85;
assign vis_psp_o[8] = M92m85;
assign J0m675 = Ab2m85;
assign vis_r0_o[11] = Pc2m85;
assign vis_r1_o[11] = Ee2m85;
assign vis_r2_o[11] = Tf2m85;
assign vis_r3_o[11] = Ih2m85;
assign vis_r8_o[11] = Xi2m85;
assign vis_r9_o[11] = Mk2m85;
assign vis_r10_o[11] = Bm2m85;
assign vis_r11_o[11] = Qn2m85;
assign vis_r4_o[11] = Fp2m85;
assign vis_r5_o[11] = Uq2m85;
assign vis_r6_o[11] = Js2m85;
assign vis_r7_o[11] = Yt2m85;
assign vis_pc_o[11] = Nv2m85;
assign vis_r12_o[11] = Zw2m85;
assign vis_r14_o[11] = Oy2m85;
assign vis_msp_o[9] = D03m85;
assign vis_psp_o[9] = R13m85;
assign Yg2l85[11] = F33m85;
assign Pf2l85[11] = V43m85;
assign V72l85[11] = M63m85;
assign U1m675 = D83m85;
assign vis_r0_o[12] = S93m85;
assign vis_r1_o[12] = Hb3m85;
assign vis_r2_o[12] = Wc3m85;
assign vis_r3_o[12] = Le3m85;
assign vis_r8_o[12] = Ag3m85;
assign vis_r9_o[12] = Ph3m85;
assign vis_r10_o[12] = Ej3m85;
assign vis_r11_o[12] = Tk3m85;
assign vis_r4_o[12] = Im3m85;
assign vis_r5_o[12] = Xn3m85;
assign vis_r6_o[12] = Mp3m85;
assign vis_r7_o[12] = Br3m85;
assign vis_pc_o[12] = Qs3m85;
assign vis_r12_o[12] = Cu3m85;
assign vis_r14_o[12] = Rv3m85;
assign vis_msp_o[10] = Gx3m85;
assign vis_psp_o[10] = Vy3m85;
assign Yg2l85[12] = K04m85;
assign Pf2l85[12] = A24m85;
assign V72l85[12] = R34m85;
assign Qj2l85[12] = I54m85;
assign Gi2l85[12] = A74m85;
assign F3m675 = S84m85;
assign vis_r0_o[13] = Ha4m85;
assign vis_r1_o[13] = Wb4m85;
assign vis_r2_o[13] = Ld4m85;
assign vis_r3_o[13] = Af4m85;
assign vis_r8_o[13] = Pg4m85;
assign vis_r9_o[13] = Ei4m85;
assign vis_r10_o[13] = Tj4m85;
assign vis_r11_o[13] = Il4m85;
assign vis_r4_o[13] = Xm4m85;
assign vis_r5_o[13] = Mo4m85;
assign vis_r6_o[13] = Bq4m85;
assign vis_r7_o[13] = Qr4m85;
assign vis_r12_o[13] = Ft4m85;
assign vis_r14_o[13] = Uu4m85;
assign vis_msp_o[11] = Jw4m85;
assign vis_psp_o[11] = Yx4m85;
assign Yg2l85[13] = Nz4m85;
assign Pf2l85[13] = D15m85;
assign V72l85[13] = U25m85;
assign Qj2l85[13] = L45m85;
assign Gi2l85[13] = D65m85;
assign Q4m675 = V75m85;
assign M7m675 = K95m85;
assign X8m675 = Za5m85;
assign Iam675 = Oc5m85;
assign Wim675 = De5m85;
assign Slm675 = Sf5m85;
assign Dnm675 = Hh5m85;
assign Oom675 = Wi5m85;
assign Zpm675 = Lk5m85;
assign Vsm675 = Am5m85;
assign Zmo675 = Pn5m85;
assign vis_r0_o[22] = Bp5m85;
assign vis_r1_o[22] = Qq5m85;
assign vis_r2_o[22] = Fs5m85;
assign vis_r3_o[22] = Ut5m85;
assign vis_r8_o[22] = Jv5m85;
assign vis_r9_o[22] = Yw5m85;
assign vis_r10_o[22] = Ny5m85;
assign vis_r11_o[22] = C06m85;
assign vis_r4_o[22] = R16m85;
assign vis_r5_o[22] = G36m85;
assign vis_r6_o[22] = V46m85;
assign vis_r7_o[22] = K66m85;
assign vis_r12_o[22] = Z76m85;
assign vis_r14_o[22] = O96m85;
assign vis_msp_o[20] = Db6m85;
assign vis_psp_o[20] = Sc6m85;
assign Agm675 = He6m85;
assign vis_r12_o[21] = Wf6m85;
assign vis_r14_o[21] = Lh6m85;
assign vis_msp_o[19] = Aj6m85;
assign vis_psp_o[19] = Pk6m85;
assign Pem675 = Em6m85;
assign vis_r12_o[20] = Tn6m85;
assign vis_r14_o[20] = Ip6m85;
assign vis_msp_o[18] = Xq6m85;
assign vis_psp_o[18] = Ms6m85;
assign Edm675 = Bu6m85;
assign vis_r12_o[19] = Qv6m85;
assign vis_r14_o[19] = Fx6m85;
assign vis_msp_o[17] = Uy6m85;
assign vis_psp_o[17] = J07m85;
assign Tbm675 = Y17m85;
assign V72l85[23] = N37m85;
assign Qj2l85[9] = E57m85;
assign Qj2l85[25] = V67m85;
assign vis_r12_o[25] = N87m85;
assign vis_r14_o[25] = Ca7m85;
assign vis_msp_o[23] = Rb7m85;
assign vis_psp_o[23] = Gd7m85;
assign Hkm675 = Ve7m85;
assign vis_r12_o[15] = Kg7m85;
assign vis_r14_o[15] = Zh7m85;
assign vis_msp_o[13] = Oj7m85;
assign vis_psp_o[13] = Dl7m85;
assign B6m675 = Sm7m85;
assign Uhp675 = Ho7m85;
assign Lhm675 = Xp7m85;
assign sys_reset_req_o = Mr7m85;
assign Wfr675 = (!Mr7m85);
assign Vc2l85 = (V72l85 - 1'b1);
assign {R32l85, Al2l85} = ({D7n675, R5n675, F4n675, T2n675, H1n675, 
 Vzm675, Jym675, Xwm675, M2s675} - 1'b1);
assign E52l85 = (vis_pc_o + 1'b1);
assign {Nx1l85, Yl2l85} = ({vis_pc_o[30:2], Hoo675} + 1'b1);
assign {Wm2l85, Un2l85, So2l85, Qp2l85, Oq2l85, Mr2l85, Ks2l85, It2l85, 
 Gu2l85, Fv2l85, Ew2l85, Dx2l85, Cy2l85, Bz2l85, A03l85, Z03l85, 
 Y13l85, X23l85, W33l85, V43l85, U53l85, T63l85, S73l85, R83l85, 
 Q93l85, Pa3l85, Ob3l85, Nc3l85, Md3l85, Le3l85, Kf3l85, Jg3l85, 
 Tz1l85} = (J22l85 * B12l85);
assign Dt7m85 = ({{I7j675, L8j675, O9j675, Raj675, Ubj675, Xcj675,
 Aej675, Dfj675, Ggj675, Jhj675, Mij675, Pjj675, Skj675, Vlj675,
 Ymj675, Boj675, Epj675, Hqj675, Krj675, Nsj675, Qtj675, Tuj675,
 Wvj675, Zwj675, Cyj675, Fzj675, I0k675, K1k675, M2k675, O3k675,
 Q4k675, S5k675, U6k675}, 1'b0} + {{1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, W7k675}, 1'b1});
assign {F6j675, Sy1l85} = Dt7m85[33:1];
assign Tu7m85 = ({{1'b0, Rjl675, Gil675, Vgl675, Kfl675, Zdl675, Ocl675,
 Dbl675, S9l675, H8l675, W6l675, L5l675, A4l675, P2l675, E1l675,
 Tzk675, Iyk675, Xwk675, Mvk675, Buk675, Qsk675, Frk675, Upk675,
 Kok675, Ank675, Qlk675, Gkk675, Wik675, Mhk675, Cgk675, Sek675,
 Idk675, Ybk675}, 1'b0} + {{1'b0, Kq1l85, Nak675, Yq1l85, Rq1l85,
 Fr1l85, As1l85, Tr1l85, Mr1l85, Os1l85, Uv1l85, Nv1l85, Bw1l85,
 Gv1l85, Zu1l85, Lu1l85, Eu1l85, Su1l85, Xt1l85, Qt1l85, Jt1l85,
 Ct1l85, Vs1l85, Pp1l85, Wp1l85, Ip1l85, Dq1l85, No1l85, Uo1l85,
 F2s675, Bp1l85, Hs1l85, D9k675}, 1'b1});
assign {I7j675, L8j675, O9j675, Raj675, Ubj675, Xcj675, Aej675, Dfj675, 
 Ggj675, Jhj675, Mij675, Pjj675, Skj675, Vlj675, Ymj675, Boj675, 
 Epj675, Hqj675, Krj675, Nsj675, Qtj675, Tuj675, Wvj675, Zwj675, 
 Cyj675, Fzj675, I0k675, K1k675, M2k675, O3k675, Q4k675, S5k675, 
 U6k675} = Tu7m85[33:1];
assign D7n675 = (Csn675 & P8n675);
assign R5n675 = (Rqn675 & P8n675);
assign F4n675 = (Gpn675 & P8n675);
assign T2n675 = (Vnn675 & P8n675);
assign H1n675 = (Lmn675 & P8n675);
assign Vzm675 = (Bln675 & P8n675);
assign Jym675 = (Rjn675 & P8n675);
assign Xwm675 = (Hin675 & P8n675);
assign Hoo675 = (~(A4y675 & H4y675));
assign H4y675 = (~(vis_pc_o[1] & O4y675));
assign B12l85[9] = (~(V4y675 | C5y675));
assign B12l85[8] = (~(C5y675 | J5y675));
assign B12l85[7] = (~(C5y675 | Q5y675));
assign B12l85[6] = (~(C5y675 | X5y675));
assign B12l85[5] = (~(C5y675 | E6y675));
assign B12l85[4] = (~(C5y675 | L6y675));
assign B12l85[3] = (~(C5y675 | S6y675));
assign B12l85[31] = (~(C5y675 | Z6y675));
assign B12l85[30] = (~(C5y675 | G7y675));
assign B12l85[2] = (~(C5y675 | N7y675));
assign B12l85[29] = (~(C5y675 | U7y675));
assign B12l85[28] = (~(C5y675 | B8y675));
assign B12l85[27] = (~(C5y675 | I8y675));
assign B12l85[26] = (~(C5y675 | P8y675));
assign B12l85[25] = (~(C5y675 | W8y675));
assign B12l85[24] = (~(C5y675 | D9y675));
assign B12l85[23] = (~(K9y675 | C5y675));
assign B12l85[22] = (~(C5y675 | R9y675));
assign B12l85[21] = (~(C5y675 | Y9y675));
assign B12l85[20] = (~(C5y675 | Fay675));
assign B12l85[1] = (~(C5y675 | May675));
assign B12l85[19] = (~(C5y675 | Tay675));
assign B12l85[18] = (~(C5y675 | Aby675));
assign B12l85[17] = (~(C5y675 | Hby675));
assign B12l85[16] = (~(C5y675 | Oby675));
assign B12l85[15] = (~(C5y675 | Vby675));
assign B12l85[14] = (~(C5y675 | Ccy675));
assign B12l85[13] = (~(C5y675 | Jcy675));
assign B12l85[12] = (~(C5y675 | Qcy675));
assign B12l85[11] = (~(C5y675 | Xcy675));
assign B12l85[10] = (~(C5y675 | Edy675));
assign B12l85[0] = (~(C5y675 | Ldy675));
assign J22l85[9] = (~(C5y675 | Sdy675));
assign J22l85[8] = (~(C5y675 | Zdy675));
assign J22l85[7] = (~(C5y675 | Gey675));
assign J22l85[6] = (~(C5y675 | Ney675));
assign J22l85[5] = (~(C5y675 | Uey675));
assign J22l85[4] = (~(C5y675 | Bfy675));
assign J22l85[3] = (~(C5y675 | Ify675));
assign J22l85[31] = (~(C5y675 | Pfy675));
assign J22l85[30] = (~(C5y675 | Wfy675));
assign J22l85[2] = (~(C5y675 | Dgy675));
assign J22l85[29] = (~(C5y675 | Kgy675));
assign J22l85[28] = (~(C5y675 | Rgy675));
assign J22l85[27] = (~(C5y675 | Ygy675));
assign J22l85[26] = (~(C5y675 | Fhy675));
assign J22l85[25] = (~(C5y675 | Mhy675));
assign J22l85[24] = (~(C5y675 | Thy675));
assign J22l85[23] = (~(C5y675 | Aiy675));
assign J22l85[22] = (~(C5y675 | Hiy675));
assign J22l85[21] = (~(C5y675 | Oiy675));
assign J22l85[20] = (~(C5y675 | Viy675));
assign J22l85[1] = (~(C5y675 | Cjy675));
assign J22l85[19] = (~(C5y675 | Jjy675));
assign J22l85[18] = (~(C5y675 | Qjy675));
assign J22l85[17] = (~(C5y675 | Xjy675));
assign J22l85[16] = (~(C5y675 | Eky675));
assign J22l85[15] = (~(C5y675 | Lky675));
assign J22l85[14] = (~(C5y675 | Sky675));
assign J22l85[13] = (~(C5y675 | Zky675));
assign J22l85[12] = (~(C5y675 | Gly675));
assign J22l85[11] = (~(C5y675 | Nly675));
assign J22l85[10] = (~(C5y675 | Uly675));
assign J22l85[0] = (~(C5y675 | Bmy675));
assign C5y675 = (Imy675 & Pmy675);
assign Pmy675 = (~(Wmy675 & Dny675));
assign Wmy675 = (Bvh675 & Kny675);
assign Imy675 = (Rny675 | Lrh675);
assign Kok675 = (~(Yny675 | Foy675));
assign Ank675 = (~(Moy675 | Foy675));
assign Qlk675 = (~(Toy675 | Foy675));
assign Gkk675 = (~(Apy675 | Foy675));
assign Wik675 = (~(Hpy675 | Foy675));
assign Mhk675 = (~(Opy675 | Foy675));
assign Cgk675 = (~(Vpy675 | Foy675));
assign Gil675 = (Cqy675 & Jqy675);
assign Sek675 = (Qqy675 & Xqy675);
assign Qqy675 = (Ery675 & Jqy675);
assign Ery675 = (~(Lry675 & Sry675));
assign Lry675 = (Gvo675 & Zry675);
assign Vgl675 = (~(Gsy675 | Foy675));
assign Kfl675 = (~(Nsy675 | Foy675));
assign Zdl675 = (~(Usy675 | Foy675));
assign Ocl675 = (~(Bty675 | Foy675));
assign Dbl675 = (~(Ity675 | Foy675));
assign S9l675 = (~(Pty675 | Foy675));
assign H8l675 = (~(Wty675 | Foy675));
assign W6l675 = (~(Duy675 | Foy675));
assign L5l675 = (~(Kuy675 | Foy675));
assign A4l675 = (~(Ruy675 | Foy675));
assign Idk675 = (~(Yuy675 | Foy675));
assign P2l675 = (~(Fvy675 | Foy675));
assign E1l675 = (~(Mvy675 | Foy675));
assign Tzk675 = (~(Tvy675 | Foy675));
assign Iyk675 = (~(Awy675 | Foy675));
assign Xwk675 = (~(Hwy675 | Foy675));
assign Mvk675 = (~(Owy675 | Foy675));
assign Buk675 = (~(Vwy675 | Foy675));
assign Qsk675 = (~(Cxy675 | Foy675));
assign Frk675 = (~(Jxy675 | Foy675));
assign Upk675 = (~(Qxy675 | Foy675));
assign Ybk675 = (~(Xxy675 | Foy675));
assign W7k675 = (Gvo675 & Eyy675);
assign Eyy675 = (~(Lyy675 & Syy675));
assign Syy675 = (Zyy675 & Gzy675);
assign Gzy675 = (~(Nzy675 & Uzy675));
assign Uzy675 = (~(B0z675 & I0z675));
assign I0z675 = (~(P0z675 & W0z675));
assign W0z675 = (~(D1z675 | K1z675));
assign P0z675 = (~(R1z675 | Y1z675));
assign Zyy675 = (~(Bvh675 & F2z675));
assign F2z675 = (~(M2z675 & T2z675));
assign T2z675 = (~(A3z675 & Mwo675));
assign M2z675 = (~(vis_apsr_o[1] & H3z675));
assign H3z675 = (~(O3z675 & V3z675));
assign V3z675 = (C4z675 | O4p675);
assign O3z675 = (Y1z675 | Ezo675);
assign Lyy675 = (J4z675 & Q4z675);
assign Q4z675 = (X4z675 | N0p675);
assign sleeping_o = (Uhp675 & E5z675);
assign T3y675 = (L5z675 ? Pf2l85[23] : hwdata_o[23]);
assign M3y675 = (~(S5z675 & Z5z675));
assign Z5z675 = (G6z675 | hready_i);
assign S5z675 = (N6z675 & U6z675);
assign N6z675 = (~(B7z675 & I7z675));
assign F3y675 = (P7z675 & irq_i[0]);
assign P7z675 = (W7z675 & D8z675);
assign D8z675 = (~(K8z675 & R8z675));
assign W7z675 = (~(Y8z675 & F9z675));
assign F9z675 = (M9z675 | T9z675);
assign Y8z675 = (Aaz675 & Haz675);
assign Aaz675 = (~(Oaz675 & Vaz675));
assign Oaz675 = (Cbz675 | Jbz675);
assign Y2y675 = (~(Qbz675 & Xbz675));
assign Xbz675 = (~(P8n675 & Ecz675));
assign Ecz675 = (Lcz675 | Scz675);
assign R2y675 = (Zcz675 | Gdz675);
assign Zcz675 = (Udz675 ? Ndz675 : Jwn675);
assign K2y675 = (Bez675 | Iez675);
assign Iez675 = (Wez675 ? Pez675 : Gwh675);
assign Pez675 = (~(Dfz675 | Kfz675));
assign Bez675 = (~(Rfz675 & Yfz675));
assign Yfz675 = (~(Eko675 & Fgz675));
assign Rfz675 = (~(Mgz675 & Jwn675));
assign D2y675 = (~(Tgz675 & Ahz675));
assign Ahz675 = (Hhz675 | hready_i);
assign Tgz675 = (Ohz675 & U6z675);
assign Ohz675 = (~(B7z675 & Vhz675));
assign Vhz675 = (haddr_o[7] | haddr_o[2]);
assign W1y675 = (~(Ciz675 & Jiz675));
assign Jiz675 = (~(Ycr675 & Lcz675));
assign Ciz675 = (Qiz675 & U6z675);
assign Qiz675 = (~(B7z675 & Xiz675));
assign Xiz675 = (haddr_o[5] | haddr_o[3]);
assign P1y675 = (~(Ejz675 & Ljz675));
assign Ljz675 = (Sjz675 | hready_i);
assign Ejz675 = (Zjz675 & U6z675);
assign Zjz675 = (~(B7z675 & Gkz675));
assign Gkz675 = (~(haddr_o[3] ^ Nkz675));
assign I1y675 = (~(Ukz675 & Blz675));
assign Blz675 = (Ilz675 | hready_i);
assign Ukz675 = (Plz675 & U6z675);
assign U6z675 = (~(B7z675 & Wlz675));
assign Wlz675 = (~(Dmz675 & Kmz675));
assign Kmz675 = (Rmz675 & Ymz675);
assign Ymz675 = (Fnz675 & Mnz675);
assign Mnz675 = (~(Tnz675 | haddr_o[25]));
assign Tnz675 = (haddr_o[16] | haddr_o[12]);
assign Fnz675 = (~(haddr_o[26] | haddr_o[27]));
assign Rmz675 = (Aoz675 & Hoz675);
assign Hoz675 = (~(haddr_o[23] | haddr_o[24]));
assign Aoz675 = (~(haddr_o[21] | haddr_o[22]));
assign Dmz675 = (Ooz675 & Voz675);
assign Voz675 = (Cpz675 & Jpz675);
assign Jpz675 = (~(Qpz675 | haddr_o[18]));
assign Qpz675 = (haddr_o[19] | haddr_o[20]);
assign Cpz675 = (~(Xpz675 | haddr_o[17]));
assign Xpz675 = (!hsize_o[1]);
assign Ooz675 = (Eqz675 & Lqz675);
assign Lqz675 = (haddr_o[14] & haddr_o[15]);
assign Eqz675 = (Sqz675 & haddr_o[13]);
assign Sqz675 = (~(Zqz675 & Grz675));
assign Grz675 = (~(Nrz675 & Urz675));
assign Urz675 = (Bsz675 & Isz675);
assign Bsz675 = (Psz675 | Wsz675);
assign Nrz675 = (Dtz675 & Ktz675);
assign Ktz675 = (~(I7z675 ^ haddr_o[9]));
assign Dtz675 = (haddr_o[11] ? Ytz675 : Rtz675);
assign Ytz675 = (Fuz675 & haddr_o[10]);
assign Rtz675 = (Muz675 & Psz675);
assign Psz675 = (Tuz675 & Avz675);
assign Tuz675 = (~(haddr_o[6] | haddr_o[2]));
assign Muz675 = (~(haddr_o[10] | haddr_o[5]));
assign Zqz675 = (Hvz675 | Ovz675);
assign Ovz675 = (I7z675 ? haddr_o[11] : Vvz675);
assign Vvz675 = (~(Cwz675 & haddr_o[10]));
assign Cwz675 = (haddr_o[2] & haddr_o[11]);
assign Hvz675 = (~(Wsz675 & Jwz675));
assign Jwz675 = (~(Qwz675 & Nkz675));
assign Qwz675 = (~(haddr_o[4] | haddr_o[3]));
assign Wsz675 = (Xwz675 & Fuz675);
assign Fuz675 = (~(haddr_o[7] | haddr_o[9]));
assign Xwz675 = (~(haddr_o[5] | haddr_o[6]));
assign Plz675 = (~(B7z675 & Avz675));
assign B1y675 = (~(Exz675 & Lxz675));
assign Lxz675 = (~(Yg2l85[31] & Sxz675));
assign Sxz675 = (~(hwdata_o[31] & Zxz675));
assign Exz675 = (Gyz675 | Nyz675);
assign U0y675 = (~(Uyz675 & Bzz675));
assign Bzz675 = (~(Yg2l85[0] & Izz675));
assign Izz675 = (~(hwdata_o[0] & Zxz675));
assign Uyz675 = (Gyz675 | Vaz675);
assign N0y675 = (~(Pzz675 & Wzz675));
assign Wzz675 = (D00775 & K00775);
assign K00775 = (~(R00775 & vis_tbit_o));
assign D00775 = (~(vis_pc_o[23] & Y00775));
assign Pzz675 = (F10775 & M10775);
assign M10775 = (~(T10775 & haddr_o[24]));
assign F10775 = (A20775 | H20775);
assign G0y675 = (V20775 ? vis_tbit_o : O20775);
assign V20775 = (C30775 & J30775);
assign J30775 = (~(Q30775 & X30775));
assign X30775 = (E40775 & L40775);
assign E40775 = (~(S40775 & Z40775));
assign Z40775 = (G50775 & N50775);
assign G50775 = (U50775 | Mwo675);
assign S40775 = (B60775 & I60775);
assign I60775 = (Y1z675 | K1z675);
assign B60775 = (Ezo675 | X5p675);
assign Q30775 = (~(P60775 | W60775));
assign C30775 = (D70775 | Lcz675);
assign O20775 = (~(K70775 & R70775));
assign R70775 = (Y70775 | F80775);
assign Y70775 = (!Sy1l85[0]);
assign K70775 = (M80775 & T80775);
assign T80775 = (A90775 | H90775);
assign M80775 = (D70775 | O90775);
assign Zzx675 = (~(V90775 & Ca0775));
assign Ca0775 = (Ja0775 & Qa0775);
assign Qa0775 = (~(Xa0775 & hrdata_i[15]));
assign Ja0775 = (Eb0775 & Lb0775);
assign Lb0775 = (~(Tio675 & Fgz675));
assign Eb0775 = (~(Sb0775 & hrdata_i[31]));
assign V90775 = (Zb0775 & Gc0775);
assign Gc0775 = (~(Yun675 & Mgz675));
assign Zb0775 = (Nc0775 | Wez675);
assign Szx675 = (~(Uc0775 & Bd0775));
assign Bd0775 = (Id0775 & Pd0775);
assign Pd0775 = (~(hrdata_i[13] & Xa0775));
assign Id0775 = (Wd0775 & De0775);
assign De0775 = (~(Xfo675 & Fgz675));
assign Wd0775 = (~(hrdata_i[29] & Sb0775));
assign Uc0775 = (Ke0775 & Re0775);
assign Re0775 = (~(Mgz675 & Csn675));
assign Ke0775 = (Ye0775 | Wez675);
assign Lzx675 = (Mf0775 ? Hsi675 : Ff0775);
assign Ff0775 = (~(Tf0775 & Ag0775));
assign Ag0775 = (Hg0775 & Og0775);
assign Og0775 = (Vg0775 & Ch0775);
assign Vg0775 = (~(Jh0775 | Sry675));
assign Hg0775 = (Qh0775 & Xh0775);
assign Xh0775 = (~(Ei0775 & Li0775));
assign Ei0775 = (Si0775 ^ Zi0775);
assign Qh0775 = (Gj0775 & Nj0775);
assign Nj0775 = (~(Uj0775 & Bk0775));
assign Uj0775 = (Ik0775 & Ye0775);
assign Gj0775 = (~(Pk0775 & Wk0775));
assign Pk0775 = (~(K1z675 | F3p675));
assign Tf0775 = (Dl0775 & Kl0775);
assign Kl0775 = (Rl0775 & Yl0775);
assign Yl0775 = (Fm0775 | Mm0775);
assign Rl0775 = (Tm0775 & An0775);
assign An0775 = (~(Z9n675 & Hn0775));
assign Tm0775 = (On0775 | Vn0775);
assign Dl0775 = (Co0775 & Jo0775);
assign Jo0775 = (~(Qo0775 & Xo0775));
assign Co0775 = (Ep0775 | W1p675);
assign Ezx675 = (Sp0775 ? vis_r0_o[1] : Lp0775);
assign Xyx675 = (Gq0775 ? Zp0775 : vis_apsr_o[1]);
assign Gq0775 = (hready_i & Nq0775);
assign Nq0775 = (~(Uq0775 & Br0775));
assign Zp0775 = (~(Ir0775 & Pr0775));
assign Pr0775 = (D70775 | Wr0775);
assign Ir0775 = (Ds0775 & Ks0775);
assign Ks0775 = (~(Br0775 & Rs0775));
assign Ds0775 = (~(Ys0775 & Ft0775));
assign Qyx675 = (~(Mt0775 & Tt0775));
assign Tt0775 = (Au0775 & Hu0775);
assign Hu0775 = (~(R00775 & vis_apsr_o[1]));
assign Au0775 = (~(Y00775 & vis_pc_o[28]));
assign Mt0775 = (Ou0775 & Vu0775);
assign Vu0775 = (~(T10775 & haddr_o[29]));
assign Ou0775 = (Cv0775 | H20775);
assign Jyx675 = (~(Jv0775 & Qv0775));
assign Qv0775 = (~(Xv0775 & Br0775));
assign Jv0775 = (hready_i ? Lw0775 : Ew0775);
assign Lw0775 = (~(Sw0775 & Zw0775));
assign Zw0775 = (~(Gx0775 & Br0775));
assign Sw0775 = (Br0775 ? Ux0775 : Nx0775);
assign Ux0775 = (By0775 & Iy0775);
assign Iy0775 = (~(Rjl675 & Sy1l85[31]));
assign By0775 = (Kq1l85 ? Rjl675 : Sy1l85[31]);
assign Nx0775 = (Py0775 & Wy0775);
assign Wy0775 = (~(Dz0775 & Kz0775));
assign Kz0775 = (D70775 | Rz0775);
assign Py0775 = (~(Rz0775 & Yz0775));
assign Ew0775 = (!vis_apsr_o[0]);
assign Cyx675 = (~(F01775 & M01775));
assign M01775 = (T01775 & A11775);
assign A11775 = (~(vis_apsr_o[0] & R00775));
assign T01775 = (~(Y00775 & vis_pc_o[27]));
assign F01775 = (H11775 & O11775);
assign O11775 = (~(T10775 & haddr_o[28]));
assign H11775 = (V11775 | H20775);
assign Vxx675 = (Sp0775 ? vis_r0_o[28] : C21775);
assign Oxx675 = (Sp0775 ? vis_r0_o[31] : J21775);
assign Hxx675 = (~(Q21775 & X21775));
assign X21775 = (E31775 | H20775);
assign Q21775 = (L31775 & S31775);
assign S31775 = (~(vis_pc_o[6] & Y00775));
assign L31775 = (~(T10775 & haddr_o[7]));
assign Axx675 = (Sp0775 ? vis_r0_o[7] : Z31775);
assign Twx675 = (Sp0775 ? vis_r0_o[0] : G41775);
assign Mwx675 = (U41775 ? N41775 : M62l85[0]);
assign N41775 = (!B51775);
assign Fwx675 = (~(I51775 & P51775));
assign P51775 = (~(W51775 & D61775));
assign D61775 = (K61775 & R61775);
assign W51775 = (U41775 & Y61775);
assign I51775 = (~(F71775 & Lcz675));
assign F71775 = (~(M71775 & T71775));
assign T71775 = (~(hresp_i & A81775));
assign A81775 = (~(H81775 & O81775));
assign O81775 = (V81775 & C91775);
assign C91775 = (~(J91775 & Q91775));
assign J91775 = (~(X91775 & Ea1775));
assign Ea1775 = (~(La1775 & Sa1775));
assign La1775 = (~(Za1775 | X5p675));
assign V81775 = (Gb1775 & Nb1775);
assign Gb1775 = (~(Ub1775 & Bc1775));
assign Bc1775 = (~(Ic1775 & Pc1775));
assign Pc1775 = (~(Wc1775 & Dd1775));
assign Dd1775 = (~(Kd1775 & Rd1775));
assign Kd1775 = (Yd1775 & Fe1775);
assign Fe1775 = (Me1775 | Ezo675);
assign Yd1775 = (Te1775 | R1z675);
assign Ic1775 = (Af1775 | Vxo675);
assign H81775 = (Hf1775 & Of1775);
assign Hf1775 = (Vf1775 & Cg1775);
assign Cg1775 = (~(O4p675 & Jg1775));
assign Jg1775 = (~(Qg1775 & Xg1775));
assign Xg1775 = (~(Eh1775 & Zry675));
assign Qg1775 = (~(Lh1775 & Sh1775));
assign Vf1775 = (Zh1775 | Af1775);
assign Yvx675 = (Gi1775 ? vis_r1_o[31] : J21775);
assign Rvx675 = (Gi1775 ? vis_r1_o[28] : C21775);
assign Kvx675 = (Gi1775 ? vis_r1_o[7] : Z31775);
assign Dvx675 = (Gi1775 ? vis_r1_o[1] : Lp0775);
assign Wux675 = (Gi1775 ? vis_r1_o[0] : G41775);
assign Pux675 = (Ui1775 ? Ni1775 : vis_primask_o);
assign Ui1775 = (~(Lcz675 | Bj1775));
assign Iux675 = (~(Ij1775 & Pj1775));
assign Pj1775 = (Wj1775 & Dk1775);
assign Dk1775 = (~(Xa0775 & hrdata_i[0]));
assign Wj1775 = (Kk1775 & Rk1775);
assign Rk1775 = (~(Uxn675 & Fgz675));
assign Kk1775 = (~(Sb0775 & hrdata_i[16]));
assign Ij1775 = (Yk1775 & Fl1775);
assign Fl1775 = (~(Z9n675 & Mgz675));
assign Yk1775 = (Fm0775 | Wez675);
assign Bux675 = (Mf0775 ? Lti675 : Ml1775);
assign Ml1775 = (~(Tl1775 & Am1775));
assign Am1775 = (Hm1775 & Om1775);
assign Om1775 = (Vm1775 & Ch0775);
assign Vm1775 = (~(Cn1775 & Li0775));
assign Cn1775 = (Jn1775 ^ Qn1775);
assign Hm1775 = (Xn1775 & Eo1775);
assign Eo1775 = (~(Lo1775 & Qo0775));
assign Lo1775 = (~(So1775 ^ Hsi675));
assign Xn1775 = (~(Jbn675 & Hn0775));
assign Tl1775 = (Zo1775 & Gp1775);
assign Gp1775 = (Np1775 & Up1775);
assign Up1775 = (~(Bq1775 & T7i675));
assign Np1775 = (Iq1775 | Vn0775);
assign Zo1775 = (Pq1775 & Wq1775);
assign Wq1775 = (Dr1775 | Mm0775);
assign Pq1775 = (~(Kr1775 & Jfi675));
assign Utx675 = (~(Rr1775 & Yr1775));
assign Yr1775 = (~(Fs1775 & hready_i));
assign Fs1775 = (Ms1775 & Ts1775);
assign Ms1775 = (~(At1775 & Ht1775));
assign Rr1775 = (E5z675 | Ot1775);
assign Ntx675 = (~(Vt1775 & Cu1775));
assign Cu1775 = (~(Ju1775 & Ts1775));
assign Vt1775 = (Qu1775 & Xu1775);
assign Xu1775 = (~(Z9n675 & Ev1775));
assign Qu1775 = (~(Lv1775 & hrdata_i[0]));
assign Gtx675 = (~(Sv1775 & Zv1775));
assign Zv1775 = (Gw1775 | Nw1775);
assign Sv1775 = (Uw1775 & Bx1775);
assign Bx1775 = (~(Ix1775 & Z9n675));
assign Uw1775 = (Px1775 | A90775);
assign Zsx675 = (~(Wx1775 & Dy1775));
assign Dy1775 = (~(Ky1775 & Ts1775));
assign Wx1775 = (Ry1775 & Yy1775);
assign Yy1775 = (~(Jbn675 & Ev1775));
assign Ry1775 = (~(Lv1775 & hrdata_i[1]));
assign Ssx675 = (~(Fz1775 & Mz1775));
assign Mz1775 = (Tz1775 | Nw1775);
assign Fz1775 = (A02775 & H02775);
assign H02775 = (~(Ix1775 & Jbn675));
assign A02775 = (Px1775 | O02775);
assign Lsx675 = (~(V02775 & C12775));
assign C12775 = (~(J12775 & Ts1775));
assign V02775 = (Q12775 & X12775);
assign X12775 = (~(Tcn675 & Ev1775));
assign Q12775 = (~(hrdata_i[2] & Lv1775));
assign Esx675 = (~(E22775 & L22775));
assign L22775 = (~(S22775 & Ts1775));
assign E22775 = (Z22775 & G32775);
assign G32775 = (~(Den675 & Ev1775));
assign Z22775 = (~(hrdata_i[3] & Lv1775));
assign Xrx675 = (~(N32775 & U32775));
assign U32775 = (~(B42775 & Ts1775));
assign N32775 = (I42775 & P42775);
assign P42775 = (~(Nfn675 & Ev1775));
assign I42775 = (~(Lv1775 & hrdata_i[4]));
assign Qrx675 = (~(W42775 & D52775));
assign D52775 = (~(K52775 & Ts1775));
assign W42775 = (R52775 & Y52775);
assign Y52775 = (~(Xgn675 & Ev1775));
assign Ev1775 = (~(Udz675 & F62775));
assign F62775 = (Ts1775 | M62775);
assign R52775 = (~(Lv1775 & hrdata_i[5]));
assign Jrx675 = (~(T62775 & A72775));
assign A72775 = (~(H72775 & Hin675));
assign T62775 = (O72775 & V72775);
assign V72775 = (~(R32l85[1] & C82775));
assign O72775 = (~(hrdata_i[6] & Lv1775));
assign Crx675 = (~(J82775 & Q82775));
assign Q82775 = (~(H72775 & Rjn675));
assign J82775 = (X82775 & E92775);
assign E92775 = (~(R32l85[2] & C82775));
assign X82775 = (~(Lv1775 & hrdata_i[7]));
assign Vqx675 = (~(L92775 & S92775));
assign S92775 = (~(H72775 & Bln675));
assign L92775 = (Z92775 & Ga2775);
assign Ga2775 = (~(R32l85[3] & C82775));
assign Z92775 = (~(Lv1775 & hrdata_i[8]));
assign Oqx675 = (~(Na2775 & Ua2775));
assign Ua2775 = (~(H72775 & Lmn675));
assign Na2775 = (Bb2775 & Ib2775);
assign Ib2775 = (~(R32l85[4] & C82775));
assign Bb2775 = (~(Lv1775 & hrdata_i[9]));
assign Hqx675 = (~(Pb2775 & Wb2775));
assign Wb2775 = (~(H72775 & Vnn675));
assign Pb2775 = (Dc2775 & Kc2775);
assign Kc2775 = (~(R32l85[5] & C82775));
assign Dc2775 = (~(hrdata_i[10] & Lv1775));
assign Aqx675 = (~(Rc2775 & Yc2775));
assign Yc2775 = (~(H72775 & Gpn675));
assign Rc2775 = (Fd2775 & Md2775);
assign Md2775 = (~(R32l85[6] & C82775));
assign Fd2775 = (~(hrdata_i[11] & Lv1775));
assign Tpx675 = (~(Td2775 & Ae2775));
assign Ae2775 = (~(H72775 & Rqn675));
assign Td2775 = (He2775 & Oe2775);
assign Oe2775 = (~(R32l85[7] & C82775));
assign He2775 = (~(Lv1775 & hrdata_i[12]));
assign Mpx675 = (~(Ve2775 & Cf2775));
assign Cf2775 = (~(H72775 & Csn675));
assign Ve2775 = (Jf2775 & Qf2775);
assign Qf2775 = (~(R32l85[8] & C82775));
assign C82775 = (Xf2775 & Gdz675);
assign Xf2775 = (~(Ts1775 & Eg2775));
assign Eg2775 = (~(Lg2775 & Sg2775));
assign Sg2775 = (Zg2775 & Gh2775);
assign Gh2775 = (P8n675 & Nh2775);
assign Nh2775 = (~(Jbn675 ^ Ky1775));
assign Zg2775 = (Uh2775 & Bi2775);
assign Bi2775 = (~(J12775 ^ Tcn675));
assign Uh2775 = (~(B42775 ^ Nfn675));
assign Lg2775 = (Ii2775 & Pi2775);
assign Pi2775 = (~(Ju1775 ^ Z9n675));
assign Ii2775 = (Wi2775 & Dj2775);
assign Dj2775 = (~(S22775 ^ Den675));
assign Wi2775 = (~(K52775 ^ Xgn675));
assign Jf2775 = (~(Lv1775 & hrdata_i[13]));
assign Fpx675 = (~(Kj2775 & Rj2775));
assign Rj2775 = (~(hrdata_i[14] & Lv1775));
assign Lv1775 = (Yj2775 & Kfz675);
assign Yj2775 = (~(Gdz675 | H72775));
assign Kj2775 = (~(Ntn675 & H72775));
assign Yox675 = (Fk2775 | Gdz675);
assign Fk2775 = (H72775 ? Yun675 : Mk2775);
assign Mk2775 = (Kfz675 & hrdata_i[15]);
assign Rox675 = (!Tk2775);
assign Tk2775 = (H72775 ? Al2775 : Gdz675);
assign H72775 = (!Udz675);
assign Udz675 = (~(M62775 & Hl2775));
assign Hl2775 = (~(Ol2775 & Vl2775));
assign Vl2775 = (O4y675 & Cm2775);
assign Ol2775 = (~(Jm2775 | Qm2775));
assign M62775 = (!Gdz675);
assign Al2775 = (~(Xm2775 & Nvm675));
assign Xm2775 = (~(Qm2775 | Mgz675));
assign Gdz675 = (Ts1775 | P8n675);
assign Kox675 = (~(En2775 & Ln2775));
assign Ln2775 = (Sn2775 & Zn2775);
assign Zn2775 = (~(hrdata_i[1] & Xa0775));
assign Sn2775 = (Go2775 & No2775);
assign No2775 = (~(Ezn675 & Fgz675));
assign Go2775 = (~(hrdata_i[17] & Sb0775));
assign En2775 = (Uo2775 & Bp2775);
assign Bp2775 = (~(Jbn675 & Mgz675));
assign Uo2775 = (Dr1775 | Wez675);
assign Dox675 = (~(Ip2775 & Pp2775));
assign Pp2775 = (Wp2775 & Dq2775);
assign Dq2775 = (~(hrdata_i[2] & Xa0775));
assign Wp2775 = (Kq2775 & Rq2775);
assign Rq2775 = (~(O0o675 & Fgz675));
assign Kq2775 = (~(hrdata_i[18] & Sb0775));
assign Ip2775 = (Yq2775 & Fr2775);
assign Fr2775 = (~(Tcn675 & Mgz675));
assign Yq2775 = (Mr2775 | Wez675);
assign Wnx675 = (~(Tr2775 & As2775));
assign As2775 = (Hs2775 & Os2775);
assign Os2775 = (~(hrdata_i[3] & Xa0775));
assign Hs2775 = (Vs2775 & Ct2775);
assign Ct2775 = (~(Y1o675 & Fgz675));
assign Vs2775 = (~(hrdata_i[19] & Sb0775));
assign Tr2775 = (Jt2775 & Qt2775);
assign Qt2775 = (~(Den675 & Mgz675));
assign Jt2775 = (Xt2775 | Wez675);
assign Pnx675 = (~(Eu2775 & Lu2775));
assign Lu2775 = (Su2775 & Zu2775);
assign Zu2775 = (~(hrdata_i[4] & Xa0775));
assign Su2775 = (Gv2775 & Nv2775);
assign Nv2775 = (~(I3o675 & Fgz675));
assign Gv2775 = (~(hrdata_i[20] & Sb0775));
assign Eu2775 = (Uv2775 & Bw2775);
assign Bw2775 = (~(Nfn675 & Mgz675));
assign Uv2775 = (Iw2775 | Wez675);
assign Inx675 = (~(Pw2775 & Ww2775));
assign Ww2775 = (Dx2775 & Kx2775);
assign Kx2775 = (~(hrdata_i[5] & Xa0775));
assign Dx2775 = (Rx2775 & Yx2775);
assign Yx2775 = (~(S4o675 & Fgz675));
assign Rx2775 = (~(hrdata_i[21] & Sb0775));
assign Pw2775 = (Fy2775 & My2775);
assign My2775 = (~(Xgn675 & Mgz675));
assign Fy2775 = (Ty2775 | Wez675);
assign Bnx675 = (~(Az2775 & Hz2775));
assign Hz2775 = (Oz2775 & Vz2775);
assign Vz2775 = (~(hrdata_i[6] & Xa0775));
assign Oz2775 = (C03775 & J03775);
assign J03775 = (~(C6o675 & Fgz675));
assign C03775 = (~(hrdata_i[22] & Sb0775));
assign Az2775 = (Q03775 & X03775);
assign X03775 = (~(Mgz675 & Hin675));
assign Q03775 = (On0775 | Wez675);
assign Umx675 = (~(E13775 & L13775));
assign L13775 = (S13775 & Z13775);
assign Z13775 = (~(Xa0775 & hrdata_i[7]));
assign S13775 = (G23775 & N23775);
assign N23775 = (~(M7o675 & Fgz675));
assign G23775 = (~(Sb0775 & hrdata_i[23]));
assign E13775 = (U23775 & B33775);
assign B33775 = (~(Mgz675 & Rjn675));
assign U23775 = (Iq1775 | Wez675);
assign Nmx675 = (~(I33775 & P33775));
assign P33775 = (W33775 & D43775);
assign D43775 = (~(Xa0775 & hrdata_i[8]));
assign W33775 = (K43775 & R43775);
assign R43775 = (~(W8o675 & Fgz675));
assign K43775 = (~(Sb0775 & hrdata_i[24]));
assign I33775 = (Y43775 & F53775);
assign F53775 = (~(Mgz675 & Bln675));
assign Y43775 = (M53775 | Wez675);
assign Gmx675 = (~(T53775 & A63775));
assign A63775 = (H63775 & O63775);
assign O63775 = (~(hrdata_i[9] & Xa0775));
assign H63775 = (V63775 & C73775);
assign C73775 = (~(Gao675 & Fgz675));
assign V63775 = (~(hrdata_i[25] & Sb0775));
assign T53775 = (J73775 & Q73775);
assign Q73775 = (~(Mgz675 & Lmn675));
assign J73775 = (X73775 | Wez675);
assign Zlx675 = (~(E83775 & L83775));
assign L83775 = (S83775 & Z83775);
assign Z83775 = (~(hrdata_i[10] & Xa0775));
assign S83775 = (G93775 & N93775);
assign N93775 = (~(Qbo675 & Fgz675));
assign G93775 = (~(hrdata_i[26] & Sb0775));
assign E83775 = (U93775 & Ba3775);
assign Ba3775 = (~(Mgz675 & Vnn675));
assign U93775 = (Ia3775 | Wez675);
assign Slx675 = (~(Pa3775 & Wa3775));
assign Wa3775 = (Db3775 & Kb3775);
assign Kb3775 = (~(hrdata_i[11] & Xa0775));
assign Db3775 = (Rb3775 & Yb3775);
assign Yb3775 = (~(Bdo675 & Fgz675));
assign Rb3775 = (~(hrdata_i[27] & Sb0775));
assign Pa3775 = (Fc3775 & Mc3775);
assign Mc3775 = (~(Mgz675 & Gpn675));
assign Fc3775 = (Tc3775 | Wez675);
assign Llx675 = (~(Ad3775 & Hd3775));
assign Hd3775 = (Od3775 & Vd3775);
assign Vd3775 = (~(hrdata_i[12] & Xa0775));
assign Od3775 = (Ce3775 & Je3775);
assign Je3775 = (~(Meo675 & Fgz675));
assign Ce3775 = (~(hrdata_i[28] & Sb0775));
assign Ad3775 = (Qe3775 & Xe3775);
assign Xe3775 = (~(Mgz675 & Rqn675));
assign Qe3775 = (Ef3775 | Wez675);
assign Elx675 = (~(Lf3775 & Sf3775));
assign Sf3775 = (Zf3775 & Gg3775);
assign Gg3775 = (~(hrdata_i[14] & Xa0775));
assign Xa0775 = (Ng3775 & Ug3775);
assign Ug3775 = (~(Dfz675 | Bh3775));
assign Ng3775 = (~(Ndz675 | Ih3775));
assign Zf3775 = (Ph3775 & Wh3775);
assign Wh3775 = (~(Iho675 & Fgz675));
assign Fgz675 = (Di3775 & Wez675);
assign Di3775 = (Ki3775 & Dfz675);
assign Dfz675 = (!Plo675);
assign Ki3775 = (~(Ri3775 & Yi3775));
assign Yi3775 = (Fj3775 | Nvm675);
assign Ph3775 = (~(hrdata_i[30] & Sb0775));
assign Sb0775 = (Mj3775 & Kfz675);
assign Mj3775 = (Bh3775 & Wez675);
assign Bh3775 = (vis_pc_o[0] & Cm2775);
assign Lf3775 = (Tj3775 & Ak3775);
assign Ak3775 = (~(Ntn675 & Mgz675));
assign Mgz675 = (Nvm675 & Wez675);
assign Tj3775 = (Hk3775 | Wez675);
assign Wez675 = (!Ih3775);
assign Ih3775 = (~(Ok3775 & Vk3775));
assign Vk3775 = (Cl3775 & Jl3775);
assign Ok3775 = (Ql3775 & Xl3775);
assign Ql3775 = (Em3775 & Lm3775);
assign Lm3775 = (~(Sm3775 & Zm3775));
assign Zm3775 = (~(Gn3775 & Nn3775));
assign Gn3775 = (~(Qm2775 | O4y675));
assign Xkx675 = (B7z675 ? hwrite_o : Un3775);
assign B7z675 = (Bo3775 & Io3775);
assign Io3775 = (Po3775 & Wo3775);
assign Wo3775 = (~(Dp3775 | haddr_o[28]));
assign Po3775 = (Xl3775 & Kp3775);
assign Bo3775 = (Rp3775 & Yp3775);
assign Rp3775 = (~(Fq3775 | Mq3775));
assign Un3775 = (Tq3775 & Ar3775);
assign Tq3775 = (~(Hr3775 | Or3775));
assign Qkx675 = (~(Vr3775 & Cs3775));
assign Cs3775 = (~(Yg2l85[30] & Js3775));
assign Js3775 = (~(hwdata_o[30] & Zxz675));
assign Vr3775 = (Gyz675 | Qs3775);
assign Jkx675 = (~(Xs3775 & Et3775));
assign Et3775 = (~(Yg2l85[29] & Lt3775));
assign Lt3775 = (~(hwdata_o[29] & Zxz675));
assign Xs3775 = (Gyz675 | St3775);
assign Ckx675 = (~(Zt3775 & Gu3775));
assign Gu3775 = (~(Yg2l85[28] & Nu3775));
assign Nu3775 = (~(hwdata_o[28] & Zxz675));
assign Zt3775 = (Gyz675 | Uu3775);
assign Vjx675 = (~(Bv3775 & Iv3775));
assign Iv3775 = (~(Yg2l85[27] & Pv3775));
assign Pv3775 = (~(hwdata_o[27] & Zxz675));
assign Bv3775 = (Gyz675 | Wv3775);
assign Ojx675 = (~(Dw3775 & Kw3775));
assign Kw3775 = (~(Yg2l85[26] & Rw3775));
assign Rw3775 = (~(hwdata_o[26] & Zxz675));
assign Dw3775 = (Gyz675 | Yw3775);
assign Hjx675 = (~(Fx3775 & Mx3775));
assign Mx3775 = (~(Yg2l85[25] & Tx3775));
assign Tx3775 = (~(hwdata_o[25] & Zxz675));
assign Fx3775 = (Gyz675 | Ay3775);
assign Ajx675 = (~(Hy3775 & Oy3775));
assign Oy3775 = (~(Yg2l85[24] & Vy3775));
assign Vy3775 = (~(hwdata_o[24] & Zxz675));
assign Hy3775 = (Gyz675 | Cz3775);
assign Tix675 = (~(Jz3775 & Qz3775));
assign Qz3775 = (~(Yg2l85[23] & Xz3775));
assign Xz3775 = (~(hwdata_o[23] & Zxz675));
assign Jz3775 = (Gyz675 | E04775);
assign Mix675 = (~(L04775 & S04775));
assign S04775 = (~(Yg2l85[22] & Z04775));
assign Z04775 = (~(hwdata_o[22] & Zxz675));
assign L04775 = (Gyz675 | G14775);
assign Fix675 = (~(N14775 & U14775));
assign U14775 = (~(Yg2l85[21] & B24775));
assign B24775 = (~(hwdata_o[21] & Zxz675));
assign N14775 = (~(I24775 & hwdata_o[21]));
assign Yhx675 = (~(P24775 & W24775));
assign W24775 = (~(Yg2l85[20] & D34775));
assign D34775 = (~(hwdata_o[20] & Zxz675));
assign P24775 = (~(I24775 & hwdata_o[20]));
assign Rhx675 = (~(K34775 & R34775));
assign R34775 = (~(Yg2l85[19] & Y34775));
assign Y34775 = (~(hwdata_o[19] & Zxz675));
assign K34775 = (~(I24775 & hwdata_o[19]));
assign Khx675 = (~(F44775 & M44775));
assign M44775 = (~(Yg2l85[18] & T44775));
assign T44775 = (~(hwdata_o[18] & Zxz675));
assign F44775 = (Gyz675 | A54775);
assign Dhx675 = (~(H54775 & O54775));
assign O54775 = (~(Yg2l85[17] & V54775));
assign V54775 = (~(hwdata_o[17] & Zxz675));
assign H54775 = (Gyz675 | C64775);
assign Wgx675 = (~(J64775 & Q64775));
assign Q64775 = (~(Yg2l85[16] & X64775));
assign X64775 = (~(hwdata_o[16] & Zxz675));
assign J64775 = (~(I24775 & hwdata_o[16]));
assign Pgx675 = (~(E74775 & L74775));
assign L74775 = (~(Yg2l85[15] & S74775));
assign S74775 = (~(hwdata_o[15] & Zxz675));
assign E74775 = (Gyz675 | Z74775);
assign Igx675 = (~(G84775 & N84775));
assign N84775 = (~(Yg2l85[14] & U84775));
assign U84775 = (~(hwdata_o[14] & Zxz675));
assign G84775 = (Gyz675 | B94775);
assign Bgx675 = (~(I94775 & P94775));
assign P94775 = (~(Yg2l85[13] & W94775));
assign W94775 = (~(hwdata_o[13] & Zxz675));
assign I94775 = (Gyz675 | Da4775);
assign Ufx675 = (~(Ka4775 & Ra4775));
assign Ra4775 = (~(Yg2l85[12] & Ya4775));
assign Ya4775 = (~(hwdata_o[12] & Zxz675));
assign Ka4775 = (Gyz675 | Fb4775);
assign Nfx675 = (~(Mb4775 & Tb4775));
assign Tb4775 = (~(Yg2l85[11] & Ac4775));
assign Ac4775 = (~(hwdata_o[11] & Zxz675));
assign Mb4775 = (Gyz675 | Hc4775);
assign Gfx675 = (~(Oc4775 & Vc4775));
assign Vc4775 = (~(Yg2l85[10] & Cd4775));
assign Cd4775 = (~(hwdata_o[10] & Zxz675));
assign Oc4775 = (Gyz675 | Jd4775);
assign Zex675 = (~(Qd4775 & Xd4775));
assign Xd4775 = (~(Yg2l85[9] & Ee4775));
assign Ee4775 = (~(hwdata_o[9] & Zxz675));
assign Qd4775 = (~(I24775 & hwdata_o[9]));
assign Sex675 = (~(Le4775 & Se4775));
assign Se4775 = (~(Yg2l85[8] & Ze4775));
assign Ze4775 = (~(hwdata_o[8] & Zxz675));
assign Le4775 = (Gyz675 | Gf4775);
assign Lex675 = (~(Nf4775 & Uf4775));
assign Uf4775 = (~(Yg2l85[7] & Bg4775));
assign Bg4775 = (~(hwdata_o[7] & Zxz675));
assign Nf4775 = (~(I24775 & hwdata_o[7]));
assign Eex675 = (~(Ig4775 & Pg4775));
assign Pg4775 = (~(Yg2l85[6] & Wg4775));
assign Wg4775 = (~(hwdata_o[6] & Zxz675));
assign Ig4775 = (~(I24775 & hwdata_o[6]));
assign Xdx675 = (~(Dh4775 & Kh4775));
assign Kh4775 = (~(Yg2l85[5] & Rh4775));
assign Rh4775 = (~(hwdata_o[5] & Zxz675));
assign Dh4775 = (Gyz675 | Yh4775);
assign Qdx675 = (~(Fi4775 & Mi4775));
assign Mi4775 = (~(Yg2l85[4] & Ti4775));
assign Ti4775 = (~(hwdata_o[4] & Zxz675));
assign Fi4775 = (Gyz675 | Aj4775);
assign Jdx675 = (~(Hj4775 & Oj4775));
assign Oj4775 = (~(Yg2l85[3] & Vj4775));
assign Vj4775 = (~(hwdata_o[3] & Zxz675));
assign Hj4775 = (~(I24775 & hwdata_o[3]));
assign Cdx675 = (~(Ck4775 & Jk4775));
assign Jk4775 = (~(Yg2l85[2] & Qk4775));
assign Qk4775 = (~(Xk4775 & Zxz675));
assign Ck4775 = (~(I24775 & Xk4775));
assign Vcx675 = (~(El4775 & Ll4775));
assign Ll4775 = (~(Yg2l85[1] & Sl4775));
assign Sl4775 = (~(hwdata_o[1] & Zxz675));
assign Zxz675 = (~(Gyz675 & Zl4775));
assign Zl4775 = (~(Gm4775 & Nm4775));
assign Gyz675 = (!I24775);
assign El4775 = (~(I24775 & hwdata_o[1]));
assign I24775 = (Um4775 & Nm4775);
assign Um4775 = (~(Bn4775 | Or3775));
assign Ocx675 = (In4775 ? S5r675 : hwdata_o[0]);
assign Hcx675 = (In4775 ? F4r675 : hwdata_o[1]);
assign Acx675 = (In4775 ? S2r675 : Xk4775);
assign In4775 = (~(Pn4775 & Lnh675));
assign Tbx675 = (L5z675 ? Pf2l85[0] : hwdata_o[0]);
assign Mbx675 = (L5z675 ? Pf2l85[1] : hwdata_o[1]);
assign Fbx675 = (L5z675 ? Pf2l85[2] : Xk4775);
assign Yax675 = (L5z675 ? Pf2l85[3] : hwdata_o[3]);
assign Rax675 = (L5z675 ? Pf2l85[4] : hwdata_o[4]);
assign Kax675 = (L5z675 ? Pf2l85[5] : hwdata_o[5]);
assign Dax675 = (L5z675 ? Pf2l85[6] : hwdata_o[6]);
assign W9x675 = (L5z675 ? Pf2l85[7] : hwdata_o[7]);
assign P9x675 = (L5z675 ? Pf2l85[8] : hwdata_o[8]);
assign I9x675 = (L5z675 ? Pf2l85[9] : hwdata_o[9]);
assign B9x675 = (L5z675 ? Pf2l85[10] : hwdata_o[10]);
assign U8x675 = (L5z675 ? Pf2l85[11] : hwdata_o[11]);
assign N8x675 = (L5z675 ? Pf2l85[12] : hwdata_o[12]);
assign G8x675 = (L5z675 ? Pf2l85[13] : hwdata_o[13]);
assign Z7x675 = (L5z675 ? Pf2l85[14] : hwdata_o[14]);
assign S7x675 = (L5z675 ? Pf2l85[15] : hwdata_o[15]);
assign L7x675 = (L5z675 ? Pf2l85[16] : hwdata_o[16]);
assign E7x675 = (L5z675 ? Pf2l85[17] : hwdata_o[17]);
assign X6x675 = (L5z675 ? Pf2l85[18] : hwdata_o[18]);
assign Q6x675 = (L5z675 ? Pf2l85[19] : hwdata_o[19]);
assign J6x675 = (L5z675 ? Pf2l85[20] : hwdata_o[20]);
assign C6x675 = (L5z675 ? Pf2l85[21] : hwdata_o[21]);
assign V5x675 = (L5z675 ? Pf2l85[22] : hwdata_o[22]);
assign L5z675 = (~(Wn4775 & Lnh675));
assign O5x675 = (~(Do4775 & Ko4775));
assign Ko4775 = (~(Ro4775 & V72l85[0]));
assign Do4775 = (Yo4775 & Fp4775);
assign Fp4775 = (~(Vc2l85[0] & Mp4775));
assign Yo4775 = (~(Tp4775 & Pf2l85[0]));
assign H5x675 = (~(Aq4775 & Hq4775));
assign Hq4775 = (~(Ro4775 & V72l85[1]));
assign Aq4775 = (Oq4775 & Vq4775);
assign Vq4775 = (~(Vc2l85[1] & Mp4775));
assign Oq4775 = (~(Tp4775 & Pf2l85[1]));
assign A5x675 = (~(Cr4775 & Jr4775));
assign Jr4775 = (~(V72l85[2] & Ro4775));
assign Cr4775 = (Qr4775 & Xr4775);
assign Xr4775 = (~(Vc2l85[2] & Mp4775));
assign Qr4775 = (~(Tp4775 & Pf2l85[2]));
assign T4x675 = (~(Es4775 & Ls4775));
assign Ls4775 = (~(V72l85[3] & Ro4775));
assign Es4775 = (Ss4775 & Zs4775);
assign Zs4775 = (~(Vc2l85[3] & Mp4775));
assign Ss4775 = (~(Tp4775 & Pf2l85[3]));
assign M4x675 = (~(Gt4775 & Nt4775));
assign Nt4775 = (~(Ro4775 & V72l85[4]));
assign Gt4775 = (Ut4775 & Bu4775);
assign Bu4775 = (~(Vc2l85[4] & Mp4775));
assign Ut4775 = (~(Tp4775 & Pf2l85[4]));
assign F4x675 = (~(Iu4775 & Pu4775));
assign Pu4775 = (~(Ro4775 & V72l85[5]));
assign Iu4775 = (Wu4775 & Dv4775);
assign Dv4775 = (~(Vc2l85[5] & Mp4775));
assign Wu4775 = (~(Tp4775 & Pf2l85[5]));
assign Y3x675 = (~(Kv4775 & Rv4775));
assign Rv4775 = (~(V72l85[6] & Ro4775));
assign Kv4775 = (Yv4775 & Fw4775);
assign Fw4775 = (~(Vc2l85[6] & Mp4775));
assign Yv4775 = (~(Tp4775 & Pf2l85[6]));
assign R3x675 = (~(Mw4775 & Tw4775));
assign Tw4775 = (~(Ro4775 & V72l85[7]));
assign Mw4775 = (Ax4775 & Hx4775);
assign Hx4775 = (~(Vc2l85[7] & Mp4775));
assign Ax4775 = (~(Tp4775 & Pf2l85[7]));
assign K3x675 = (~(Ox4775 & Vx4775));
assign Vx4775 = (~(Ro4775 & V72l85[8]));
assign Ox4775 = (Cy4775 & Jy4775);
assign Jy4775 = (~(Vc2l85[8] & Mp4775));
assign Cy4775 = (~(Tp4775 & Pf2l85[8]));
assign D3x675 = (~(Qy4775 & Xy4775));
assign Xy4775 = (~(Ro4775 & V72l85[9]));
assign Qy4775 = (Ez4775 & Lz4775);
assign Lz4775 = (~(Vc2l85[9] & Mp4775));
assign Ez4775 = (~(Tp4775 & Pf2l85[9]));
assign W2x675 = (~(Sz4775 & Zz4775));
assign Zz4775 = (~(V72l85[10] & Ro4775));
assign Sz4775 = (G05775 & N05775);
assign N05775 = (~(Vc2l85[10] & Mp4775));
assign G05775 = (~(Tp4775 & Pf2l85[10]));
assign P2x675 = (~(U05775 & B15775));
assign B15775 = (~(V72l85[11] & Ro4775));
assign U05775 = (I15775 & P15775);
assign P15775 = (~(Vc2l85[11] & Mp4775));
assign I15775 = (~(Tp4775 & Pf2l85[11]));
assign I2x675 = (~(W15775 & D25775));
assign D25775 = (~(Ro4775 & V72l85[12]));
assign W15775 = (K25775 & R25775);
assign R25775 = (~(Vc2l85[12] & Mp4775));
assign K25775 = (~(Tp4775 & Pf2l85[12]));
assign B2x675 = (~(Y25775 & F35775));
assign F35775 = (~(Ro4775 & V72l85[13]));
assign Y25775 = (M35775 & T35775);
assign T35775 = (~(Vc2l85[13] & Mp4775));
assign M35775 = (~(Tp4775 & Pf2l85[13]));
assign U1x675 = (~(A45775 & H45775));
assign H45775 = (~(V72l85[14] & Ro4775));
assign A45775 = (O45775 & V45775);
assign V45775 = (~(Vc2l85[14] & Mp4775));
assign O45775 = (~(Tp4775 & Pf2l85[14]));
assign N1x675 = (~(C55775 & J55775));
assign J55775 = (~(Ro4775 & V72l85[15]));
assign C55775 = (Q55775 & X55775);
assign X55775 = (~(Vc2l85[15] & Mp4775));
assign Q55775 = (~(Tp4775 & Pf2l85[15]));
assign G1x675 = (~(E65775 & L65775));
assign L65775 = (~(Ro4775 & V72l85[16]));
assign E65775 = (S65775 & Z65775);
assign Z65775 = (~(Vc2l85[16] & Mp4775));
assign S65775 = (~(Tp4775 & Pf2l85[16]));
assign Z0x675 = (~(G75775 & N75775));
assign N75775 = (~(Ro4775 & V72l85[17]));
assign G75775 = (U75775 & B85775);
assign B85775 = (~(Vc2l85[17] & Mp4775));
assign U75775 = (~(Tp4775 & Pf2l85[17]));
assign S0x675 = (~(I85775 & P85775));
assign P85775 = (~(V72l85[18] & Ro4775));
assign I85775 = (W85775 & D95775);
assign D95775 = (~(Vc2l85[18] & Mp4775));
assign W85775 = (~(Tp4775 & Pf2l85[18]));
assign L0x675 = (~(K95775 & R95775));
assign R95775 = (~(V72l85[19] & Ro4775));
assign K95775 = (Y95775 & Fa5775);
assign Fa5775 = (~(Vc2l85[19] & Mp4775));
assign Y95775 = (~(Tp4775 & Pf2l85[19]));
assign E0x675 = (~(Ma5775 & Ta5775));
assign Ta5775 = (~(Ro4775 & V72l85[20]));
assign Ma5775 = (Ab5775 & Hb5775);
assign Hb5775 = (~(Vc2l85[20] & Mp4775));
assign Ab5775 = (~(Tp4775 & Pf2l85[20]));
assign Xzw675 = (~(Ob5775 & Vb5775));
assign Vb5775 = (~(Ro4775 & V72l85[21]));
assign Ob5775 = (Cc5775 & Jc5775);
assign Jc5775 = (~(Vc2l85[21] & Mp4775));
assign Cc5775 = (~(Tp4775 & Pf2l85[21]));
assign Qzw675 = (~(Qc5775 & Xc5775));
assign Xc5775 = (~(V72l85[22] & Ro4775));
assign Qc5775 = (Ed5775 & Ld5775);
assign Ld5775 = (~(Vc2l85[22] & Mp4775));
assign Ed5775 = (~(Tp4775 & Pf2l85[22]));
assign Jzw675 = (~(Sd5775 & Zd5775));
assign Zd5775 = (~(Ro4775 & V72l85[23]));
assign Sd5775 = (Ge5775 & Ne5775);
assign Ne5775 = (~(Vc2l85[23] & Mp4775));
assign Mp4775 = (~(Ue5775 | Bf5775));
assign Ue5775 = (Ro4775 | If5775);
assign Ge5775 = (~(Tp4775 & Pf2l85[23]));
assign Tp4775 = (Pf5775 & Bf5775);
assign Bf5775 = (~(Wf5775 | V72l85[0]));
assign Pf5775 = (~(Ro4775 | If5775));
assign Ro4775 = (~(Dg5775 | If5775));
assign Czw675 = (Kg5775 ? Mb2l85[56] : hwdata_o[6]);
assign Vyw675 = (Kg5775 ? Mb2l85[57] : hwdata_o[7]);
assign Oyw675 = (Kg5775 ? Mb2l85[58] : hwdata_o[14]);
assign Hyw675 = (Kg5775 ? Mb2l85[59] : hwdata_o[15]);
assign Ayw675 = (Kg5775 ? Mb2l85[60] : hwdata_o[22]);
assign Txw675 = (Kg5775 ? Mb2l85[61] : hwdata_o[23]);
assign Mxw675 = (Kg5775 ? Mb2l85[62] : hwdata_o[30]);
assign Fxw675 = (Kg5775 ? Mb2l85[63] : hwdata_o[31]);
assign Kg5775 = (~(Rg5775 & Lnh675));
assign Yww675 = (Yg5775 ? Mb2l85[48] : hwdata_o[6]);
assign Rww675 = (Yg5775 ? Mb2l85[49] : hwdata_o[7]);
assign Kww675 = (Yg5775 ? Mb2l85[50] : hwdata_o[14]);
assign Dww675 = (Yg5775 ? Mb2l85[51] : hwdata_o[15]);
assign Wvw675 = (Yg5775 ? Mb2l85[52] : hwdata_o[22]);
assign Pvw675 = (Yg5775 ? Mb2l85[53] : hwdata_o[23]);
assign Ivw675 = (Yg5775 ? Mb2l85[54] : hwdata_o[30]);
assign Bvw675 = (Yg5775 ? Mb2l85[55] : hwdata_o[31]);
assign Yg5775 = (~(Fh5775 & Lnh675));
assign Uuw675 = (Mh5775 ? Mb2l85[40] : hwdata_o[6]);
assign Nuw675 = (Mh5775 ? Mb2l85[41] : hwdata_o[7]);
assign Guw675 = (Mh5775 ? Mb2l85[42] : hwdata_o[14]);
assign Ztw675 = (Mh5775 ? Mb2l85[43] : hwdata_o[15]);
assign Stw675 = (Mh5775 ? Mb2l85[44] : hwdata_o[22]);
assign Ltw675 = (Mh5775 ? Mb2l85[45] : hwdata_o[23]);
assign Etw675 = (Mh5775 ? Mb2l85[46] : hwdata_o[30]);
assign Xsw675 = (Mh5775 ? Mb2l85[47] : hwdata_o[31]);
assign Mh5775 = (~(Th5775 & Lnh675));
assign Qsw675 = (Ai5775 ? Mb2l85[32] : hwdata_o[6]);
assign Jsw675 = (Ai5775 ? Mb2l85[33] : hwdata_o[7]);
assign Csw675 = (Ai5775 ? Mb2l85[34] : hwdata_o[14]);
assign Vrw675 = (Ai5775 ? Mb2l85[35] : hwdata_o[15]);
assign Orw675 = (Ai5775 ? Mb2l85[36] : hwdata_o[22]);
assign Hrw675 = (Ai5775 ? Mb2l85[37] : hwdata_o[23]);
assign Arw675 = (Ai5775 ? Mb2l85[38] : hwdata_o[30]);
assign Tqw675 = (Ai5775 ? Mb2l85[39] : hwdata_o[31]);
assign Ai5775 = (~(Hi5775 & Lnh675));
assign Mqw675 = (Oi5775 ? Mb2l85[24] : hwdata_o[6]);
assign Fqw675 = (Oi5775 ? Mb2l85[25] : hwdata_o[7]);
assign Ypw675 = (Oi5775 ? Mb2l85[26] : hwdata_o[14]);
assign Rpw675 = (Oi5775 ? Mb2l85[27] : hwdata_o[15]);
assign Kpw675 = (Oi5775 ? Mb2l85[28] : hwdata_o[22]);
assign Dpw675 = (Oi5775 ? Mb2l85[29] : hwdata_o[23]);
assign Wow675 = (Oi5775 ? Mb2l85[30] : hwdata_o[30]);
assign Pow675 = (Oi5775 ? Mb2l85[31] : hwdata_o[31]);
assign Oi5775 = (~(Vi5775 & Lnh675));
assign Iow675 = (Cj5775 ? Mb2l85[16] : hwdata_o[6]);
assign Bow675 = (Cj5775 ? Mb2l85[17] : hwdata_o[7]);
assign Unw675 = (Cj5775 ? Mb2l85[18] : hwdata_o[14]);
assign Nnw675 = (Cj5775 ? Mb2l85[19] : hwdata_o[15]);
assign Gnw675 = (Cj5775 ? Mb2l85[20] : hwdata_o[22]);
assign Zmw675 = (Cj5775 ? Mb2l85[21] : hwdata_o[23]);
assign Smw675 = (Cj5775 ? Mb2l85[22] : hwdata_o[30]);
assign Lmw675 = (Cj5775 ? Mb2l85[23] : hwdata_o[31]);
assign Cj5775 = (~(Jj5775 & Lnh675));
assign Emw675 = (Qj5775 ? Mb2l85[8] : hwdata_o[6]);
assign Xlw675 = (Qj5775 ? Mb2l85[9] : hwdata_o[7]);
assign Qlw675 = (Qj5775 ? Mb2l85[10] : hwdata_o[14]);
assign Jlw675 = (Qj5775 ? Mb2l85[11] : hwdata_o[15]);
assign Clw675 = (Qj5775 ? Mb2l85[12] : hwdata_o[22]);
assign Vkw675 = (Qj5775 ? Mb2l85[13] : hwdata_o[23]);
assign Okw675 = (Qj5775 ? Mb2l85[14] : hwdata_o[30]);
assign Hkw675 = (Qj5775 ? Mb2l85[15] : hwdata_o[31]);
assign Qj5775 = (~(Xj5775 & Lnh675));
assign Akw675 = (Ek5775 ? Mb2l85[0] : hwdata_o[6]);
assign Tjw675 = (Ek5775 ? Mb2l85[1] : hwdata_o[7]);
assign Mjw675 = (Ek5775 ? Mb2l85[2] : hwdata_o[14]);
assign Fjw675 = (Ek5775 ? Mb2l85[3] : hwdata_o[15]);
assign Yiw675 = (Ek5775 ? Mb2l85[4] : hwdata_o[22]);
assign Riw675 = (Ek5775 ? Mb2l85[5] : hwdata_o[23]);
assign Kiw675 = (Ek5775 ? Mb2l85[6] : hwdata_o[30]);
assign Diw675 = (Ek5775 ? Mb2l85[7] : hwdata_o[31]);
assign Ek5775 = (~(Lk5775 & Lnh675));
assign Whw675 = (Sk5775 ? Nbp675 : hwdata_o[4]);
assign Phw675 = (Sk5775 ? Fap675 : Xk4775);
assign Ihw675 = (Sk5775 ? Doh675 : hwdata_o[1]);
assign Sk5775 = (~(Zk5775 & Lnh675));
assign Bhw675 = (Gl5775 ? hwdata_o[30] : Ha2l85[0]);
assign Ugw675 = (Gl5775 ? hwdata_o[31] : Ha2l85[1]);
assign Gl5775 = (Nl5775 & Lnh675);
assign Ngw675 = (Ul5775 ? C92l85[0] : hwdata_o[22]);
assign Ggw675 = (Ul5775 ? C92l85[1] : hwdata_o[23]);
assign Zfw675 = (Ul5775 ? Ge2l85[0] : hwdata_o[30]);
assign Sfw675 = (Ul5775 ? Ge2l85[1] : hwdata_o[31]);
assign Ul5775 = (~(Bm5775 & Lnh675));
assign Lfw675 = (~(Im5775 & Pm5775));
assign Pm5775 = (~(Wm5775 & I1r675));
assign Wm5775 = (~(Dn5775 | If5775));
assign If5775 = (Kn5775 & Lnh675);
assign Dn5775 = (Pn4775 & Or3775);
assign Im5775 = (~(Rn5775 & Dg5775));
assign Rn5775 = (Yn5775 & V72l85[0]);
assign Efw675 = (Fo5775 & irq_i[31]);
assign Fo5775 = (Mo5775 & To5775);
assign To5775 = (~(Ap5775 & Hp5775));
assign Mo5775 = (~(Op5775 & Vp5775));
assign Vp5775 = (M9z675 | Cq5775);
assign Op5775 = (Jq5775 & Haz675);
assign Jq5775 = (~(Qq5775 & Nyz675));
assign Qq5775 = (Cbz675 | Xq5775);
assign Xew675 = (Er5775 & irq_i[29]);
assign Er5775 = (Lr5775 & Sr5775);
assign Sr5775 = (~(Zr5775 & Gs5775));
assign Lr5775 = (~(Ns5775 & Us5775));
assign Us5775 = (Bt5775 | hwdata_o[29]);
assign Ns5775 = (It5775 & Haz675);
assign It5775 = (~(Pt5775 & Wt5775));
assign Qew675 = (~(Du5775 & Ku5775));
assign Ku5775 = (Ru5775 | Nw1775);
assign Du5775 = (Yu5775 & Fv5775);
assign Fv5775 = (~(Xgn675 & Ix1775));
assign Yu5775 = (Px1775 | Mv5775);
assign Jew675 = (Tv5775 & irq_i[19]);
assign Tv5775 = (Aw5775 & Hw5775);
assign Hw5775 = (~(Ow5775 & Vw5775));
assign Aw5775 = (~(Cx5775 & Jx5775));
assign Jx5775 = (hwdata_o[19] | Bt5775);
assign Cx5775 = (Qx5775 & Haz675);
assign Qx5775 = (~(Xx5775 & Ey5775));
assign Cew675 = (Ly5775 & irq_i[18]);
assign Ly5775 = (Sy5775 & Zy5775);
assign Zy5775 = (~(Gz5775 & Nz5775));
assign Sy5775 = (~(Uz5775 & B06775));
assign B06775 = (I06775 | M9z675);
assign Uz5775 = (P06775 & Haz675);
assign P06775 = (~(A54775 & W06775));
assign W06775 = (Cbz675 | D16775);
assign Vdw675 = (~(K16775 & R16775));
assign R16775 = (Y16775 | Nw1775);
assign K16775 = (F26775 & M26775);
assign M26775 = (~(Tcn675 & Ix1775));
assign F26775 = (Px1775 | T26775);
assign Odw675 = (A36775 & irq_i[23]);
assign A36775 = (H36775 & O36775);
assign O36775 = (~(V36775 & C46775));
assign H36775 = (~(J46775 & Q46775));
assign Q46775 = (hwdata_o[23] | Bt5775);
assign J46775 = (X46775 & Haz675);
assign X46775 = (~(E56775 & L56775));
assign Hdw675 = (S56775 & irq_i[22]);
assign S56775 = (Z56775 & G66775);
assign G66775 = (~(N66775 & U66775));
assign Z56775 = (~(B76775 & I76775));
assign I76775 = (M9z675 | P76775);
assign B76775 = (W76775 & Haz675);
assign W76775 = (~(G14775 & D86775));
assign D86775 = (Cbz675 | K86775);
assign Adw675 = (R86775 & irq_i[21]);
assign R86775 = (Y86775 & F96775);
assign F96775 = (~(M96775 & T96775));
assign Y86775 = (~(Aa6775 & Ha6775));
assign Ha6775 = (hwdata_o[21] | Bt5775);
assign Aa6775 = (Oa6775 & Haz675);
assign Oa6775 = (~(Va6775 & Cb6775));
assign Tcw675 = (Jb6775 & irq_i[20]);
assign Jb6775 = (Qb6775 & Xb6775);
assign Xb6775 = (~(Ec6775 & Lc6775));
assign Qb6775 = (~(Sc6775 & Zc6775));
assign Zc6775 = (hwdata_o[20] | Bt5775);
assign Sc6775 = (Gd6775 & Haz675);
assign Gd6775 = (~(Nd6775 & Ud6775));
assign Mcw675 = (~(Be6775 & Ie6775));
assign Ie6775 = (~(Pe6775 & hwdata_o[28]));
assign Be6775 = (~(We6775 & Ifp675));
assign We6775 = (Df6775 & Kf6775);
assign Kf6775 = (~(Pe6775 & hwdata_o[27]));
assign Df6775 = (~(Rf6775 & Yf6775));
assign Fcw675 = (~(Fg6775 & Mg6775));
assign Mg6775 = (Tg6775 | Nw1775);
assign Fg6775 = (Ah6775 & Hh6775);
assign Hh6775 = (~(Nfn675 & Ix1775));
assign Ah6775 = (Px1775 | Oh6775);
assign Ybw675 = (Vh6775 & irq_i[7]);
assign Vh6775 = (Ci6775 & Ji6775);
assign Ji6775 = (~(Qi6775 & Xi6775));
assign Ci6775 = (~(Ej6775 & Lj6775));
assign Lj6775 = (M9z675 | Sj6775);
assign Ej6775 = (Zj6775 & Haz675);
assign Zj6775 = (Gk6775 | hwdata_o[7]);
assign Gk6775 = (Bt5775 & Sj6775);
assign Rbw675 = (Nk6775 & irq_i[6]);
assign Nk6775 = (Uk6775 & Bl6775);
assign Bl6775 = (~(Il6775 & Pl6775));
assign Uk6775 = (~(Wl6775 & Dm6775));
assign Dm6775 = (Km6775 | M9z675);
assign Wl6775 = (Rm6775 & Haz675);
assign Rm6775 = (Ym6775 | hwdata_o[6]);
assign Ym6775 = (Bt5775 & Km6775);
assign Kbw675 = (Fn6775 & irq_i[5]);
assign Fn6775 = (Mn6775 & Tn6775);
assign Tn6775 = (~(Ao6775 & Ho6775));
assign Mn6775 = (~(Oo6775 & Vo6775));
assign Vo6775 = (M9z675 | Cp6775);
assign Oo6775 = (Jp6775 & Haz675);
assign Jp6775 = (~(Qp6775 & Yh4775));
assign Qp6775 = (Cbz675 | Xp6775);
assign Dbw675 = (Eq6775 & irq_i[4]);
assign Eq6775 = (Lq6775 & Sq6775);
assign Sq6775 = (~(Zq6775 & Gr6775));
assign Lq6775 = (~(Nr6775 & Ur6775));
assign Ur6775 = (Bs6775 | M9z675);
assign Nr6775 = (Is6775 & Haz675);
assign Is6775 = (~(Ps6775 & Aj4775));
assign Ps6775 = (Cbz675 | Ws6775);
assign Waw675 = (Dt6775 & irq_i[3]);
assign Dt6775 = (Kt6775 & Rt6775);
assign Rt6775 = (~(Yt6775 & Fu6775));
assign Kt6775 = (~(Mu6775 & Tu6775));
assign Tu6775 = (M9z675 | Av6775);
assign Mu6775 = (Hv6775 & Haz675);
assign Hv6775 = (Ov6775 | hwdata_o[3]);
assign Ov6775 = (Bt5775 & Av6775);
assign Paw675 = (~(Vv6775 & Cw6775));
assign Cw6775 = (Jw6775 | Nw1775);
assign Vv6775 = (Qw6775 & Xw6775);
assign Xw6775 = (~(Den675 & Ix1775));
assign Ix1775 = (Ot1775 & P8n675);
assign Ot1775 = (Nw1775 & Ht1775);
assign Ht1775 = (Ex6775 | Lx6775);
assign Qw6775 = (Px1775 | Sx6775);
assign Px1775 = (~(Nw1775 & Zx6775));
assign Iaw675 = (Gy6775 & Ny6775);
assign Ny6775 = (Uy6775 & Bz6775);
assign Uy6775 = (~(Iz6775 & Pz6775));
assign Gy6775 = (nmi_i & Wz6775);
assign Wz6775 = (Cbz675 | D07775);
assign Baw675 = (~(K07775 & R07775));
assign R07775 = (Y07775 | F17775);
assign F17775 = (Oxh675 ? T17775 : M17775);
assign M17775 = (At1775 | D07775);
assign Y07775 = (~(A27775 & V8p675));
assign K07775 = (~(Tth675 & Sm3775));
assign U9w675 = (~(H27775 & O27775));
assign O27775 = (~(Cep675 & V27775));
assign V27775 = (~(C37775 & Yf6775));
assign N9w675 = (J37775 & irq_i[15]);
assign J37775 = (Q37775 & X37775);
assign X37775 = (~(E47775 & L47775));
assign Q37775 = (~(S47775 & Z47775));
assign Z47775 = (M9z675 | G57775);
assign S47775 = (N57775 & Haz675);
assign N57775 = (~(Z74775 & U57775));
assign U57775 = (Cbz675 | B67775);
assign G9w675 = (I67775 & irq_i[14]);
assign I67775 = (P67775 & W67775);
assign W67775 = (~(D77775 & K77775));
assign P67775 = (~(R77775 & Y77775));
assign Y77775 = (F87775 | M9z675);
assign R77775 = (M87775 & Haz675);
assign M87775 = (~(B94775 & T87775));
assign T87775 = (~(Bt5775 & F87775));
assign Z8w675 = (A97775 & irq_i[13]);
assign A97775 = (H97775 & O97775);
assign O97775 = (~(V97775 & Ca7775));
assign H97775 = (~(Ja7775 & Qa7775));
assign Qa7775 = (M9z675 | Xa7775);
assign Ja7775 = (Eb7775 & Haz675);
assign Eb7775 = (~(Lb7775 & Da4775));
assign Lb7775 = (Cbz675 | Sb7775);
assign S8w675 = (Zb7775 & irq_i[12]);
assign Zb7775 = (Gc7775 & Nc7775);
assign Nc7775 = (~(Uc7775 & Bd7775));
assign Gc7775 = (~(Id7775 & Pd7775));
assign Pd7775 = (M9z675 | Wd7775);
assign Id7775 = (De7775 & Haz675);
assign De7775 = (~(Ke7775 & Fb4775));
assign Ke7775 = (Cbz675 | Re7775);
assign L8w675 = (Ye7775 & irq_i[11]);
assign Ye7775 = (Ff7775 & Mf7775);
assign Mf7775 = (~(Tf7775 & Ag7775));
assign Ff7775 = (~(Hg7775 & Og7775));
assign Og7775 = (M9z675 | Vg7775);
assign Hg7775 = (Ch7775 & Haz675);
assign Ch7775 = (~(Hc4775 & Jh7775));
assign Jh7775 = (Cbz675 | Qh7775);
assign E8w675 = (Xh7775 & irq_i[10]);
assign Xh7775 = (Ei7775 & Li7775);
assign Li7775 = (~(Si7775 & Zi7775));
assign Ei7775 = (~(Gj7775 & Nj7775));
assign Nj7775 = (M9z675 | Uj7775);
assign Gj7775 = (Bk7775 & Haz675);
assign Bk7775 = (~(Ik7775 & Jd4775));
assign Ik7775 = (Cbz675 | Pk7775);
assign X7w675 = (Wk7775 & irq_i[9]);
assign Wk7775 = (Dl7775 & Kl7775);
assign Kl7775 = (~(Rl7775 & Yl7775));
assign Dl7775 = (~(Fm7775 & Mm7775));
assign Mm7775 = (M9z675 | Tm7775);
assign Fm7775 = (An7775 & Haz675);
assign An7775 = (hwdata_o[9] | Hn7775);
assign Hn7775 = (Bt5775 & Tm7775);
assign Q7w675 = (On7775 & irq_i[8]);
assign On7775 = (Vn7775 & Co7775);
assign Co7775 = (~(Jo7775 & Qo7775));
assign Vn7775 = (~(Xo7775 & Ep7775));
assign Ep7775 = (M9z675 | Lp7775);
assign Xo7775 = (Sp7775 & Haz675);
assign Sp7775 = (~(Gf4775 & Zp7775));
assign Zp7775 = (Cbz675 | Gq7775);
assign J7w675 = (Nq7775 & irq_i[28]);
assign Nq7775 = (Uq7775 & Br7775);
assign Br7775 = (~(Ir7775 & Pr7775));
assign Uq7775 = (~(Wr7775 & Ds7775));
assign Ds7775 = (Bt5775 | hwdata_o[28]);
assign Wr7775 = (Ks7775 & Haz675);
assign Ks7775 = (~(Rs7775 & Ys7775));
assign C7w675 = (Ft7775 & irq_i[27]);
assign Ft7775 = (Mt7775 & Tt7775);
assign Tt7775 = (~(Au7775 & Hu7775));
assign Mt7775 = (~(Ou7775 & Vu7775));
assign Vu7775 = (M9z675 | Cv7775);
assign Ou7775 = (Jv7775 & Haz675);
assign Jv7775 = (~(Qv7775 & Wv3775));
assign Qv7775 = (Cbz675 | Xv7775);
assign V6w675 = (Ew7775 & irq_i[26]);
assign Ew7775 = (Lw7775 & Sw7775);
assign Sw7775 = (~(Zw7775 & Gx7775));
assign Lw7775 = (~(Nx7775 & Ux7775));
assign Ux7775 = (Bt5775 | hwdata_o[26]);
assign Nx7775 = (By7775 & Haz675);
assign By7775 = (~(Iy7775 & Py7775));
assign O6w675 = (Wy7775 & irq_i[25]);
assign Wy7775 = (Dz7775 & Kz7775);
assign Kz7775 = (~(Rz7775 & Yz7775));
assign Dz7775 = (~(F08775 & M08775));
assign M08775 = (M9z675 | T08775);
assign F08775 = (A18775 & Haz675);
assign A18775 = (~(H18775 & Ay3775));
assign H18775 = (Cbz675 | O18775);
assign H6w675 = (V18775 & irq_i[24]);
assign V18775 = (C28775 & J28775);
assign J28775 = (~(Q28775 & X28775));
assign C28775 = (~(E38775 & L38775));
assign L38775 = (Bt5775 | hwdata_o[24]);
assign E38775 = (S38775 & Haz675);
assign S38775 = (~(Z38775 & G48775));
assign A6w675 = (~(N48775 & U48775));
assign U48775 = (~(Ogp675 & B58775));
assign B58775 = (~(I58775 & Yf6775));
assign N48775 = (~(P58775 & W58775));
assign W58775 = (!D68775);
assign T5w675 = (K68775 & irq_i[2]);
assign K68775 = (R68775 & Y68775);
assign Y68775 = (~(F78775 & M78775));
assign R68775 = (~(T78775 & A88775));
assign A88775 = (Bt5775 | Xk4775);
assign T78775 = (H88775 & Haz675);
assign H88775 = (~(O88775 & V88775));
assign M5w675 = (C98775 & irq_i[1]);
assign C98775 = (J98775 & Q98775);
assign Q98775 = (~(X98775 & Ea8775));
assign J98775 = (~(La8775 & Sa8775));
assign Sa8775 = (M9z675 | Za8775);
assign La8775 = (Gb8775 & Haz675);
assign Gb8775 = (Nb8775 | hwdata_o[1]);
assign Nb8775 = (Bt5775 & Za8775);
assign F5w675 = (~(Ub8775 & Bc8775));
assign Bc8775 = (~(Ic8775 & E7r675));
assign Ic8775 = (Pc8775 & Wc8775);
assign Wc8775 = (~(Pe6775 & hwdata_o[25]));
assign Pc8775 = (~(Dd8775 & Yf6775));
assign Y4w675 = (~(Kd8775 & Rd8775));
assign Rd8775 = (~(Yd8775 & V8p675));
assign Yd8775 = (Fe8775 & Me8775);
assign Fe8775 = (~(Te8775 & Af8775));
assign Af8775 = (~(Hf8775 & C37775));
assign Hf8775 = (A27775 & Of8775);
assign Te8775 = (~(Vf8775 & Nw1775));
assign Nw1775 = (hready_i & At1775);
assign Vf8775 = (~(Cg8775 | vis_pc_o[1]));
assign Kd8775 = (~(Lsh675 & Sm3775));
assign Sm3775 = (~(hready_i & Bvh675));
assign R4w675 = (Jg8775 & irq_i[17]);
assign Jg8775 = (Qg8775 & Xg8775);
assign Xg8775 = (~(Eh8775 & Lh8775));
assign Qg8775 = (~(Sh8775 & Zh8775));
assign Zh8775 = (hwdata_o[17] | Bt5775);
assign Sh8775 = (Gi8775 & Haz675);
assign Gi8775 = (~(Ni8775 & Ui8775));
assign K4w675 = (Bj8775 & irq_i[16]);
assign Bj8775 = (Ij8775 & Pj8775);
assign Pj8775 = (~(Wj8775 & Dk8775));
assign Ij8775 = (~(Kk8775 & Rk8775));
assign Rk8775 = (Yk8775 | M9z675);
assign Kk8775 = (Fl8775 & Haz675);
assign Fl8775 = (hwdata_o[16] | Ml8775);
assign Ml8775 = (Bt5775 & Yk8775);
assign D4w675 = (Tl8775 & irq_i[30]);
assign Tl8775 = (Am8775 & Hm8775);
assign Hm8775 = (~(Om8775 & Vm8775));
assign Am8775 = (~(Cn8775 & Jn8775));
assign Jn8775 = (M9z675 | Qn8775);
assign Cn8775 = (Xn8775 & Haz675);
assign Haz675 = (M9z675 | Bt5775);
assign Xn8775 = (~(Eo8775 & Qs3775));
assign Eo8775 = (Cbz675 | Lo8775);
assign W3w675 = (~(So8775 & Zo8775));
assign Zo8775 = (Gp8775 & Np8775);
assign Np8775 = (~(T10775 & haddr_o[2]));
assign haddr_o[2] = (~(Up8775 & Bq8775));
assign Bq8775 = (~(Iq8775 & Xqy675));
assign Up8775 = (Pq8775 & Wq8775);
assign Wq8775 = (~(Dr8775 & Dp3775));
assign Dr8775 = (Kr8775 & A4y675);
assign A4y675 = (~(Rr8775 & vis_pc_o[0]));
assign Rr8775 = (~(Qm2775 | Yr8775));
assign Kr8775 = (~(Yr8775 & Fs8775));
assign Fs8775 = (Fj3775 | Qm2775);
assign Yr8775 = (~(O4y675 ^ vis_pc_o[1]));
assign Pq8775 = (~(Sy1l85[2] & Ms8775));
assign Gp8775 = (~(R00775 & vis_ipsr_o[2]));
assign So8775 = (Ts8775 & At8775);
assign At8775 = (~(Y00775 & vis_pc_o[1]));
assign Ts8775 = (~(Wnl675 & Ht8775));
assign P3w675 = (~(Ot8775 & Vt8775));
assign Vt8775 = (~(Cll675 & Ht8775));
assign Ot8775 = (Cu8775 & Ju8775);
assign Ju8775 = (~(T10775 & Qu8775));
assign Qu8775 = (~(B51775 & Xu8775));
assign Xu8775 = (~(vis_tbit_o & Ev8775));
assign Ev8775 = (Lv8775 | Sv8775);
assign Sv8775 = (Zv8775 & Gw8775);
assign Zv8775 = (~(X73775 | M53775));
assign Cu8775 = (~(R00775 & vis_ipsr_o[0]));
assign I3w675 = (~(Nw8775 & Uw8775));
assign Nw8775 = (Px8775 ? Ix8775 : Bx8775);
assign Ix8775 = (Wx8775 & Dy8775);
assign Dy8775 = (Ky8775 | Iq1775);
assign Wx8775 = (Ry8775 & Yy8775);
assign Yy8775 = (~(T7i675 & Fz8775));
assign Ry8775 = (~(Xhi675 & Mz8775));
assign B3w675 = (~(Tz8775 & A09775));
assign A09775 = (~(Px8775 & H09775));
assign H09775 = (~(O09775 & V09775));
assign V09775 = (Ky8775 | M53775);
assign O09775 = (C19775 & J19775);
assign J19775 = (~(A9i675 & Fz8775));
assign C19775 = (~(Eji675 & Mz8775));
assign Tz8775 = (Q19775 & Uw8775);
assign Q19775 = (~(R2j675 & X19775));
assign X19775 = (~(Px8775 & E29775));
assign E29775 = (Bx8775 | L29775);
assign U2w675 = (~(S29775 & Z29775));
assign Z29775 = (G39775 & Uw8775);
assign G39775 = (~(V3j675 & N39775));
assign N39775 = (~(Px8775 & U39775));
assign U39775 = (B49775 | L29775);
assign S29775 = (I49775 & P49775);
assign P49775 = (~(Px8775 & W49775));
assign W49775 = (~(D59775 & K59775));
assign K59775 = (Ky8775 | X73775);
assign D59775 = (R59775 & Y59775);
assign Y59775 = (~(Hai675 & Fz8775));
assign Fz8775 = (~(F69775 & M69775));
assign M69775 = (T69775 & A79775);
assign A79775 = (~(H79775 & O79775));
assign H79775 = (V79775 & E5z675);
assign V79775 = (C89775 | Lv8775);
assign T69775 = (~(J89775 & Q89775));
assign J89775 = (~(Ef3775 | Lki675));
assign F69775 = (X89775 & E99775);
assign R59775 = (~(Lki675 & Mz8775));
assign Mz8775 = (~(L99775 & S99775));
assign S99775 = (Z99775 & Ga9775);
assign L99775 = (Na9775 & Ua9775);
assign Ua9775 = (~(Bb9775 & Ib9775));
assign Bb9775 = (~(Pb9775 | Lrh675));
assign Na9775 = (~(Q89775 & Wb9775));
assign Wb9775 = (Ef3775 | Dc9775);
assign I49775 = (Kc9775 | L29775);
assign N2w675 = (~(Rc9775 & Yc9775));
assign Yc9775 = (Px8775 ? Md9775 : Fd9775);
assign Md9775 = (Td9775 & Ae9775);
assign Ae9775 = (He9775 & Oe9775);
assign Oe9775 = (~(Ve9775 & Dc9775));
assign He9775 = (Z99775 | Tc3775);
assign Z99775 = (~(Cf9775 & E5z675));
assign Cf9775 = (Jf9775 | Qf9775);
assign Td9775 = (Xf9775 & Eg9775);
assign Eg9775 = (Xt2775 | X89775);
assign X89775 = (Lg9775 & Sg9775);
assign Lg9775 = (~(Ve9775 & Zg9775));
assign Zg9775 = (Gh9775 & Nh9775);
assign Gh9775 = (Tc3775 | X73775);
assign Ve9775 = (Q89775 & Bni675);
assign Xf9775 = (Ky8775 | Ia3775);
assign Rc9775 = (Uh9775 & Uw8775);
assign Uw8775 = (~(Px8775 & Bi9775));
assign Bi9775 = (~(Ii9775 & Pi9775));
assign Ii9775 = (Wi9775 & Dj9775);
assign Wi9775 = (~(Kj9775 & Ik0775));
assign Kj9775 = (Rj9775 & Qgi675);
assign Px8775 = (hready_i & Yj9775);
assign Yj9775 = (~(Fk9775 & Mk9775));
assign Mk9775 = (Tk9775 & Al9775);
assign Al9775 = (Hl9775 & Ol9775);
assign Ol9775 = (Vl9775 & Cm9775);
assign Hl9775 = (Jm9775 & Qm9775);
assign Tk9775 = (Xm9775 & En9775);
assign En9775 = (Ln9775 | Sn9775);
assign Xm9775 = (Zn9775 & Go9775);
assign Go9775 = (~(No9775 & Uo9775));
assign No9775 = (Bp9775 & M53775);
assign Bp9775 = (~(Nh9775 & Ip9775));
assign Ip9775 = (~(Pp9775 & Lki675));
assign Pp9775 = (~(Wp9775 | Ty2775));
assign Zn9775 = (~(Dq9775 & Kq9775));
assign Dq9775 = (~(Cm2775 | Zqi675));
assign Fk9775 = (Rq9775 & Yq9775);
assign Yq9775 = (Fr9775 & Mr9775);
assign Mr9775 = (Tr9775 & As9775);
assign As9775 = (~(Hs9775 & Gwh675));
assign Tr9775 = (~(Os9775 & Vs9775));
assign Fr9775 = (Ct9775 & Jt9775);
assign Jt9775 = (Qt9775 | Hk3775);
assign Rq9775 = (Xt9775 & Eu9775);
assign Xt9775 = (~(Lu9775 | Su9775));
assign Lu9775 = (!Zu9775);
assign Uh9775 = (Gv9775 | L29775);
assign L29775 = (Nv9775 & Uv9775);
assign Uv9775 = (Cg8775 | U50775);
assign Nv9775 = (Bw9775 & Iw9775);
assign Bw9775 = (~(Wk0775 & Pw9775));
assign G2w675 = (Mf0775 ? Pui675 : Ww9775);
assign Ww9775 = (~(Dx9775 & Kx9775));
assign Kx9775 = (Rx9775 & Yx9775);
assign Yx9775 = (Fy9775 & Ch0775);
assign Ch0775 = (~(My9775 & Ty9775));
assign Ty9775 = (~(Az9775 & Za1775));
assign Az9775 = (Mr2775 | W1p675);
assign Fy9775 = (~(Hz9775 & Li0775));
assign Hz9775 = (Oz9775 ^ Vz9775);
assign Rx9775 = (C0a775 & J0a775);
assign J0a775 = (~(Q0a775 & Qo0775));
assign Q0a775 = (~(X0a775 ^ E1a775));
assign C0a775 = (~(Tcn675 & Hn0775));
assign Dx9775 = (L1a775 & S1a775);
assign S1a775 = (Z1a775 & G2a775);
assign G2a775 = (~(Bq1775 & A9i675));
assign Z1a775 = (M53775 | Vn0775);
assign Vn0775 = (~(N2a775 | U2a775));
assign L1a775 = (B3a775 & I3a775);
assign I3a775 = (Mr2775 | Mm0775);
assign B3a775 = (~(Kr1775 & Qgi675));
assign Z1w675 = (Mf0775 ? Tvi675 : P3a775);
assign Mf0775 = (~(hready_i & W3a775));
assign W3a775 = (~(D4a775 & K4a775));
assign K4a775 = (R4a775 & Y4a775);
assign Y4a775 = (F5a775 & M5a775);
assign M5a775 = (~(T5a775 & A6a775));
assign A6a775 = (~(E5z675 & H6a775));
assign H6a775 = (Cg8775 | O6a775);
assign F5a775 = (V6a775 & C7a775);
assign V6a775 = (~(J7a775 & Q7a775));
assign J7a775 = (~(X7a775 | Mwo675));
assign R4a775 = (E8a775 & L8a775);
assign L8a775 = (~(S8a775 & Z8a775));
assign E8a775 = (Jm9775 | Ia3775);
assign Jm9775 = (~(G9a775 & N9a775));
assign G9a775 = (~(Gwh675 | Rpi675));
assign D4a775 = (U9a775 & Baa775);
assign Baa775 = (Iaa775 & Paa775);
assign Paa775 = (~(Waa775 & Dba775));
assign Iaa775 = (Kba775 | Rba775);
assign U9a775 = (Yba775 & Fca775);
assign P3a775 = (~(Mca775 & Tca775));
assign Tca775 = (Ada775 & Hda775);
assign Hda775 = (Oda775 & Vda775);
assign Vda775 = (~(Cea775 & Qo0775));
assign Qo0775 = (~(Jea775 & Qea775));
assign Jea775 = (Xea775 & Efa775);
assign Efa775 = (~(Lfa775 & Sfa775));
assign Xea775 = (~(Wk0775 & Zfa775));
assign Cea775 = (~(Gga775 ^ Nga775));
assign Nga775 = (E1a775 & Pui675);
assign E1a775 = (~(So1775 | Xo0775));
assign Oda775 = (Uga775 & Dj9775);
assign Uga775 = (~(Bha775 & Li0775));
assign Li0775 = (~(Iha775 & Pha775));
assign Pha775 = (~(Wha775 & Dia775));
assign Wha775 = (Ik0775 & Zqi675);
assign Iha775 = (~(Kia775 & Ria775));
assign Kia775 = (Q89775 & Lki675);
assign Bha775 = (~(Yia775 & Fja775));
assign Fja775 = (Vz9775 | Oz9775);
assign Oz9775 = (~(Mja775 ^ Tja775));
assign Vz9775 = (~(Qn1775 & Jn1775));
assign Jn1775 = (~(Tja775 | Aka775));
assign Aka775 = (~(Hka775 | Oka775));
assign Qn1775 = (~(Si0775 | Zi0775));
assign Zi0775 = (~(Vka775 ^ Qgi675));
assign Yia775 = (~(Tja775 & Mja775));
assign Mja775 = (~(Cla775 & Jla775));
assign Jla775 = (Qla775 & Xla775);
assign Xla775 = (~(Ema775 & Lma775));
assign Qla775 = (Sma775 | Zma775);
assign Cla775 = (Gna775 & Nna775);
assign Nna775 = (~(Una775 & Boa775));
assign Gna775 = (Ioa775 | Poa775);
assign Tja775 = (Oka775 & Hka775);
assign Hka775 = (Lma775 ^ Ema775);
assign Ema775 = (~(On0775 | Woa775));
assign Lma775 = (Boa775 ^ Una775);
assign Una775 = (Dpa775 & Cei675);
assign Boa775 = (Poa775 ^ Ioa775);
assign Poa775 = (~(Sma775 ^ Zma775));
assign Zma775 = (~(Kpa775 | Rpa775));
assign Oka775 = (Qgi675 & Vka775);
assign Vka775 = (Woa775 ^ On0775);
assign Woa775 = (Dpa775 ^ Ty2775);
assign Dpa775 = (Ioa775 & Ypa775);
assign Ypa775 = (~(Fqa775 & Iw2775));
assign Ioa775 = (Fqa775 | Iw2775);
assign Fqa775 = (~(Sma775 & Mqa775));
assign Mqa775 = (Tqa775 | Obi675);
assign Sma775 = (~(Tqa775 & Obi675));
assign Tqa775 = (~(Kpa775 | Ara775));
assign Ara775 = (~(Hra775 | Hai675));
assign Kpa775 = (Hra775 & Hai675);
assign Hra775 = (~(Rpa775 | Ora775));
assign Ada775 = (Vra775 & Csa775);
assign Csa775 = (~(Den675 & Hn0775));
assign Hn0775 = (P8n675 & Jsa775);
assign Jsa775 = (~(Qsa775 & Xsa775));
assign Xsa775 = (Eta775 | Zfa775);
assign Vra775 = (~(Bq1775 & Hai675));
assign Bq1775 = (Ik0775 & Lta775);
assign Lta775 = (Sta775 | Uo9775);
assign Mca775 = (Zta775 & Gua775);
assign Gua775 = (Nua775 & Uua775);
assign Uua775 = (~(Eji675 & N2a775));
assign N2a775 = (~(Bva775 & Iva775));
assign Iva775 = (~(Pva775 & Nc0775));
assign Pva775 = (~(Wva775 & E99775));
assign E99775 = (Pb9775 | Dwa775);
assign Bva775 = (~(U2a775 & Tc3775));
assign Nua775 = (Xt2775 | Mm0775);
assign Mm0775 = (Kwa775 & Rwa775);
assign Rwa775 = (Ywa775 & Ga9775);
assign Ywa775 = (~(Fxa775 & Mxa775));
assign Mxa775 = (~(Tc3775 | Zqi675));
assign Fxa775 = (Ik0775 & N9a775);
assign Kwa775 = (Txa775 & Aya775);
assign Aya775 = (~(Q89775 & Hya775));
assign Hya775 = (~(Ria775 & Lki675));
assign Txa775 = (Oya775 | Vya775);
assign Zta775 = (Cza775 & Jza775);
assign Jza775 = (~(Kr1775 & Xhi675));
assign Cza775 = (~(Qza775 & Xza775));
assign S1w675 = (L0b775 ? E0i675 : E0b775);
assign E0b775 = (~(S0b775 & Z0b775));
assign Z0b775 = (G1b775 & N1b775);
assign N1b775 = (U1b775 & B2b775);
assign U1b775 = (~(I2b775 & A9i675));
assign G1b775 = (P2b775 & W2b775);
assign W2b775 = (~(D3b775 & K3b775));
assign K3b775 = (~(R3b775 & Y3b775));
assign R3b775 = (T4b775 ? M4b775 : F4b775);
assign M4b775 = (~(Bx8775 & B49775));
assign P2b775 = (~(Vci675 & A5b775));
assign S0b775 = (H5b775 & O5b775);
assign H5b775 = (V5b775 & C6b775);
assign C6b775 = (J6b775 | Iq1775);
assign V5b775 = (B49775 | Q6b775);
assign L1w675 = (X6b775 ? vis_r2_o[31] : J21775);
assign E1w675 = (X6b775 ? vis_r2_o[28] : C21775);
assign X0w675 = (X6b775 ? vis_r2_o[7] : Z31775);
assign Q0w675 = (X6b775 ? vis_r2_o[1] : Lp0775);
assign J0w675 = (X6b775 ? vis_r2_o[0] : G41775);
assign C0w675 = (E7b775 ? vis_r3_o[31] : J21775);
assign Vzv675 = (E7b775 ? vis_r3_o[28] : C21775);
assign Ozv675 = (E7b775 ? vis_r3_o[7] : Z31775);
assign Hzv675 = (E7b775 ? vis_r3_o[1] : Lp0775);
assign Azv675 = (E7b775 ? vis_r3_o[0] : G41775);
assign Tyv675 = (L7b775 ? vis_r8_o[31] : J21775);
assign Myv675 = (L7b775 ? vis_r8_o[28] : C21775);
assign Fyv675 = (L7b775 ? vis_r8_o[7] : Z31775);
assign Yxv675 = (L7b775 ? vis_r8_o[1] : Lp0775);
assign Rxv675 = (L7b775 ? vis_r8_o[0] : G41775);
assign Kxv675 = (S7b775 ? vis_r9_o[31] : J21775);
assign Dxv675 = (S7b775 ? vis_r9_o[28] : C21775);
assign Wwv675 = (S7b775 ? vis_r9_o[7] : Z31775);
assign Pwv675 = (S7b775 ? vis_r9_o[1] : Lp0775);
assign Iwv675 = (S7b775 ? vis_r9_o[0] : G41775);
assign Bwv675 = (Z7b775 ? vis_r10_o[31] : J21775);
assign Uvv675 = (Z7b775 ? vis_r10_o[28] : C21775);
assign Nvv675 = (Z7b775 ? vis_r10_o[7] : Z31775);
assign Gvv675 = (Z7b775 ? vis_r10_o[1] : Lp0775);
assign Zuv675 = (Z7b775 ? vis_r10_o[0] : G41775);
assign Suv675 = (G8b775 ? vis_r11_o[31] : J21775);
assign Luv675 = (G8b775 ? vis_r11_o[28] : C21775);
assign Euv675 = (G8b775 ? vis_r11_o[7] : Z31775);
assign Xtv675 = (G8b775 ? vis_r11_o[1] : Lp0775);
assign Qtv675 = (G8b775 ? vis_r11_o[0] : G41775);
assign Jtv675 = (N8b775 ? vis_r14_o[31] : J21775);
assign Ctv675 = (N8b775 ? vis_r14_o[28] : C21775);
assign Vsv675 = (N8b775 ? vis_r14_o[7] : Z31775);
assign Osv675 = (N8b775 ? vis_r14_o[1] : Lp0775);
assign Hsv675 = (N8b775 ? vis_r14_o[0] : G41775);
assign Asv675 = (U8b775 ? vis_r12_o[31] : J21775);
assign Trv675 = (U8b775 ? vis_r12_o[28] : C21775);
assign Mrv675 = (U8b775 ? vis_r12_o[7] : Z31775);
assign Frv675 = (U8b775 ? vis_r12_o[1] : Lp0775);
assign Yqv675 = (U8b775 ? vis_r12_o[0] : G41775);
assign Rqv675 = (B9b775 ? vis_r7_o[31] : J21775);
assign Kqv675 = (B9b775 ? vis_r7_o[28] : C21775);
assign Dqv675 = (B9b775 ? vis_r7_o[7] : Z31775);
assign Wpv675 = (B9b775 ? vis_r7_o[1] : Lp0775);
assign Ppv675 = (B9b775 ? vis_r7_o[0] : G41775);
assign Ipv675 = (I9b775 ? vis_r6_o[31] : J21775);
assign Bpv675 = (I9b775 ? vis_r6_o[28] : C21775);
assign Uov675 = (I9b775 ? vis_r6_o[7] : Z31775);
assign Nov675 = (I9b775 ? vis_r6_o[1] : Lp0775);
assign Gov675 = (I9b775 ? vis_r6_o[0] : G41775);
assign Znv675 = (P9b775 ? vis_r5_o[31] : J21775);
assign Snv675 = (P9b775 ? vis_r5_o[28] : C21775);
assign Lnv675 = (P9b775 ? vis_r5_o[7] : Z31775);
assign Env675 = (P9b775 ? vis_r5_o[1] : Lp0775);
assign Xmv675 = (P9b775 ? vis_r5_o[0] : G41775);
assign Qmv675 = (W9b775 ? vis_r4_o[31] : J21775);
assign Jmv675 = (W9b775 ? vis_r4_o[28] : C21775);
assign Cmv675 = (W9b775 ? vis_r4_o[7] : Z31775);
assign Vlv675 = (W9b775 ? vis_r4_o[1] : Lp0775);
assign Lp0775 = (~(O02775 & Dab775));
assign Olv675 = (W9b775 ? vis_r4_o[0] : G41775);
assign G41775 = (~(Kab775 & Rab775));
assign Rab775 = (Yab775 & Fbb775);
assign Fbb775 = (~(Mbb775 & Sy1l85[0]));
assign Yab775 = (Tbb775 & Acb775);
assign Acb775 = (~(Hcb775 & D9k675));
assign Hcb775 = (~(Ocb775 | Vcb775));
assign Tbb775 = (Cdb775 | Jdb775);
assign Kab775 = (A90775 & Qdb775);
assign A90775 = (Xdb775 & Eeb775);
assign Eeb775 = (Leb775 & Seb775);
assign Seb775 = (Zeb775 | Gfb775);
assign Leb775 = (Nfb775 & Ufb775);
assign Nfb775 = (Bgb775 | Igb775);
assign Xdb775 = (Pgb775 & Wgb775);
assign Wgb775 = (Dhb775 | Khb775);
assign Pgb775 = (Rhb775 | Yhb775);
assign Hlv675 = (~(Fib775 & Mib775));
assign Mib775 = (Tib775 & Ajb775);
assign Ajb775 = (~(Hjb775 & Ojb775));
assign Ojb775 = (~(Vjb775 | Ckb775));
assign Hjb775 = (~(Jkb775 | Dia775));
assign Tib775 = (~(R00775 & vis_ipsr_o[1]));
assign Fib775 = (Qkb775 & Xkb775);
assign Xkb775 = (~(Y00775 & vis_pc_o[0]));
assign Qkb775 = (Elb775 | H20775);
assign Alv675 = (Slb775 ? Llb775 : vis_control_o);
assign Slb775 = (hready_i & Zlb775);
assign Zlb775 = (~(Gmb775 & Nmb775));
assign Nmb775 = (~(Umb775 & Bnb775));
assign Bnb775 = (Xwi675 & Inb775);
assign Umb775 = (~(Pnb775 | X0a775));
assign Gmb775 = (~(Yf6775 | Wnb775));
assign Llb775 = (~(Dob775 & Kob775));
assign Kob775 = (~(Inb775 & Rob775));
assign Dob775 = (~(G5i675 & vis_pc_o[1]));
assign Tkv675 = (Fpb775 ? Yob775 : Gum675);
assign Fpb775 = (hready_i & Mpb775);
assign Mpb775 = (~(Tpb775 & Aqb775));
assign Aqb775 = (Hqb775 & Oqb775);
assign Oqb775 = (Vqb775 & Crb775);
assign Vqb775 = (Jrb775 & Qrb775);
assign Hqb775 = (Xrb775 & Esb775);
assign Esb775 = (~(Lsb775 & Ssb775));
assign Lsb775 = (Sa1775 & Kny675);
assign Xrb775 = (~(Zsb775 & Gtb775));
assign Tpb775 = (Ntb775 & Utb775);
assign Utb775 = (Bub775 & Iub775);
assign Iub775 = (Pub775 | X5p675);
assign Bub775 = (Wub775 | Xt2775);
assign Ntb775 = (Dvb775 & Kvb775);
assign Kvb775 = (~(Qza775 & Nzy675));
assign Dvb775 = (~(Rvb775 & Yvb775));
assign Yob775 = (~(Fwb775 & Mwb775));
assign Mwb775 = (~(Twb775 & Axb775));
assign Axb775 = (Hxb775 | Oxb775);
assign Oxb775 = (Ezo675 ? Vxb775 : My9775);
assign Vxb775 = (Cg8775 | Ora775);
assign Hxb775 = (~(Cyb775 & Dj9775));
assign Cyb775 = (Y1z675 ? Obi675 : W1p675);
assign Twb775 = (vis_control_o | Jyb775);
assign Jyb775 = (Wnb775 & vis_pc_o[1]);
assign Fwb775 = (T7i675 ? Xyb775 : Qyb775);
assign Xyb775 = (Vya775 | Ezo675);
assign Qyb775 = (~(Ezb775 & Lzb775));
assign Ezb775 = (~(Dr1775 | Xt2775));
assign Mkv675 = (Szb775 ? Z31775 : vis_psp_o[5]);
assign Fkv675 = (Szb775 ? C21775 : vis_psp_o[26]);
assign Yjv675 = (Szb775 ? J21775 : vis_psp_o[29]);
assign Rjv675 = (Zzb775 ? Z31775 : vis_msp_o[5]);
assign Z31775 = (~(G0c775 & N0c775));
assign Kjv675 = (Zzb775 ? C21775 : vis_msp_o[26]);
assign C21775 = (~(U0c775 & Rz0775));
assign Djv675 = (Zzb775 ? J21775 : vis_msp_o[29]);
assign J21775 = (~(B1c775 & I1c775));
assign Wiv675 = (Szb775 ? P1c775 : vis_psp_o[28]);
assign Piv675 = (Zzb775 ? P1c775 : vis_msp_o[28]);
assign Iiv675 = (N8b775 ? vis_r14_o[30] : P1c775);
assign Biv675 = (U8b775 ? vis_r12_o[30] : P1c775);
assign Uhv675 = (B9b775 ? vis_r7_o[30] : P1c775);
assign Nhv675 = (I9b775 ? vis_r6_o[30] : P1c775);
assign Ghv675 = (P9b775 ? vis_r5_o[30] : P1c775);
assign Zgv675 = (W9b775 ? vis_r4_o[30] : P1c775);
assign Sgv675 = (G8b775 ? vis_r11_o[30] : P1c775);
assign Lgv675 = (Z7b775 ? vis_r10_o[30] : P1c775);
assign Egv675 = (S7b775 ? vis_r9_o[30] : P1c775);
assign Xfv675 = (L7b775 ? vis_r8_o[30] : P1c775);
assign Qfv675 = (E7b775 ? vis_r3_o[30] : P1c775);
assign Jfv675 = (X6b775 ? vis_r2_o[30] : P1c775);
assign Cfv675 = (Gi1775 ? vis_r1_o[30] : P1c775);
assign Vev675 = (Sp0775 ? vis_r0_o[30] : P1c775);
assign P1c775 = (~(W1c775 & D2c775));
assign D2c775 = (K2c775 & R2c775);
assign R2c775 = (Cdb775 | Y2c775);
assign K2c775 = (F3c775 & M3c775);
assign F3c775 = (T3c775 | Ocb775);
assign W1c775 = (A4c775 & H4c775);
assign A4c775 = (O4c775 & V4c775);
assign V4c775 = (~(Mbb775 & Sy1l85[30]));
assign Oev675 = (J5c775 ? C5c775 : vis_apsr_o[2]);
assign C5c775 = (~(Q5c775 & X5c775));
assign X5c775 = (D70775 | H4c775);
assign Q5c775 = (E6c775 & L6c775);
assign L6c775 = (~(Br0775 & S6c775));
assign E6c775 = (Yz0775 | Y2c775);
assign Hev675 = (~(Z6c775 & G7c775));
assign G7c775 = (N7c775 & U7c775);
assign U7c775 = (~(vis_apsr_o[2] & R00775));
assign N7c775 = (~(Y00775 & vis_pc_o[29]));
assign Z6c775 = (B8c775 & I8c775);
assign I8c775 = (Jkb775 | P8c775);
assign B8c775 = (~(Krm675 & Ht8775));
assign Aev675 = (Szb775 ? W8c775 : vis_psp_o[27]);
assign Tdv675 = (Zzb775 ? W8c775 : vis_msp_o[27]);
assign Mdv675 = (N8b775 ? vis_r14_o[29] : W8c775);
assign Fdv675 = (U8b775 ? vis_r12_o[29] : W8c775);
assign Ycv675 = (B9b775 ? vis_r7_o[29] : W8c775);
assign Rcv675 = (I9b775 ? vis_r6_o[29] : W8c775);
assign Kcv675 = (P9b775 ? vis_r5_o[29] : W8c775);
assign Dcv675 = (W9b775 ? vis_r4_o[29] : W8c775);
assign Wbv675 = (G8b775 ? vis_r11_o[29] : W8c775);
assign Pbv675 = (Z7b775 ? vis_r10_o[29] : W8c775);
assign Ibv675 = (S7b775 ? vis_r9_o[29] : W8c775);
assign Bbv675 = (L7b775 ? vis_r8_o[29] : W8c775);
assign Uav675 = (E7b775 ? vis_r3_o[29] : W8c775);
assign Nav675 = (X6b775 ? vis_r2_o[29] : W8c775);
assign Gav675 = (Gi1775 ? vis_r1_o[29] : W8c775);
assign Z9v675 = (Sp0775 ? vis_r0_o[29] : W8c775);
assign W8c775 = (~(Wr0775 & D9c775));
assign S9v675 = (~(K9c775 & R9c775));
assign R9c775 = (Y9c775 | H20775);
assign K9c775 = (Fac775 & Mac775);
assign Mac775 = (~(vis_pc_o[26] & Y00775));
assign Fac775 = (~(T10775 & haddr_o[27]));
assign L9v675 = (Szb775 ? Tac775 : vis_psp_o[25]);
assign E9v675 = (Zzb775 ? Tac775 : vis_msp_o[25]);
assign X8v675 = (N8b775 ? vis_r14_o[27] : Tac775);
assign Q8v675 = (U8b775 ? vis_r12_o[27] : Tac775);
assign J8v675 = (B9b775 ? vis_r7_o[27] : Tac775);
assign C8v675 = (I9b775 ? vis_r6_o[27] : Tac775);
assign V7v675 = (P9b775 ? vis_r5_o[27] : Tac775);
assign O7v675 = (W9b775 ? vis_r4_o[27] : Tac775);
assign H7v675 = (G8b775 ? vis_r11_o[27] : Tac775);
assign A7v675 = (Z7b775 ? vis_r10_o[27] : Tac775);
assign T6v675 = (S7b775 ? vis_r9_o[27] : Tac775);
assign M6v675 = (L7b775 ? vis_r8_o[27] : Tac775);
assign F6v675 = (E7b775 ? vis_r3_o[27] : Tac775);
assign Y5v675 = (X6b775 ? vis_r2_o[27] : Tac775);
assign R5v675 = (Gi1775 ? vis_r1_o[27] : Tac775);
assign K5v675 = (Sp0775 ? vis_r0_o[27] : Tac775);
assign Tac775 = (Abc775 | Hbc775);
assign D5v675 = (~(Obc775 & Vbc775));
assign Vbc775 = (Ccc775 | H20775);
assign Obc775 = (Jcc775 & Qcc775);
assign Qcc775 = (~(vis_pc_o[25] & Y00775));
assign Jcc775 = (~(T10775 & haddr_o[26]));
assign W4v675 = (Szb775 ? Xcc775 : vis_psp_o[24]);
assign P4v675 = (Zzb775 ? Xcc775 : vis_msp_o[24]);
assign I4v675 = (N8b775 ? vis_r14_o[26] : Xcc775);
assign B4v675 = (U8b775 ? vis_r12_o[26] : Xcc775);
assign U3v675 = (B9b775 ? vis_r7_o[26] : Xcc775);
assign N3v675 = (I9b775 ? vis_r6_o[26] : Xcc775);
assign G3v675 = (P9b775 ? vis_r5_o[26] : Xcc775);
assign Z2v675 = (W9b775 ? vis_r4_o[26] : Xcc775);
assign S2v675 = (G8b775 ? vis_r11_o[26] : Xcc775);
assign L2v675 = (Z7b775 ? vis_r10_o[26] : Xcc775);
assign E2v675 = (S7b775 ? vis_r9_o[26] : Xcc775);
assign X1v675 = (L7b775 ? vis_r8_o[26] : Xcc775);
assign Q1v675 = (E7b775 ? vis_r3_o[26] : Xcc775);
assign J1v675 = (X6b775 ? vis_r2_o[26] : Xcc775);
assign C1v675 = (Gi1775 ? vis_r1_o[26] : Xcc775);
assign V0v675 = (Sp0775 ? vis_r0_o[26] : Xcc775);
assign Xcc775 = (~(Edc775 & Ldc775));
assign Ldc775 = (Sdc775 & Zdc775);
assign Zdc775 = (~(Gec775 | Tz1l85[26]));
assign Sdc775 = (Nec775 & Uec775);
assign Nec775 = (~(Bfc775 & Bty675));
assign Bfc775 = (As1l85 & Ifc775);
assign Edc775 = (Pfc775 & Wfc775);
assign Pfc775 = (Dgc775 & Kgc775);
assign Kgc775 = (Cdb775 | Rgc775);
assign Dgc775 = (~(Mbb775 & Sy1l85[26]));
assign O0v675 = (~(Ygc775 & Fhc775));
assign Fhc775 = (Mhc775 | H20775);
assign Ygc775 = (Thc775 & Aic775);
assign Aic775 = (~(vis_pc_o[24] & Y00775));
assign Thc775 = (~(T10775 & haddr_o[25]));
assign haddr_o[25] = (~(Hic775 & Oic775));
assign Oic775 = (~(Nx1l85[24] & Dp3775));
assign Hic775 = (Vic775 & Cjc775);
assign Cjc775 = (Jjc775 | Ity675);
assign Vic775 = (~(Sy1l85[25] & Ms8775));
assign H0v675 = (Szb775 ? Qjc775 : vis_psp_o[23]);
assign A0v675 = (Zzb775 ? Qjc775 : vis_msp_o[23]);
assign Tzu675 = (N8b775 ? vis_r14_o[25] : Qjc775);
assign Mzu675 = (U8b775 ? vis_r12_o[25] : Qjc775);
assign Fzu675 = (B9b775 ? vis_r7_o[25] : Qjc775);
assign Yyu675 = (I9b775 ? vis_r6_o[25] : Qjc775);
assign Ryu675 = (P9b775 ? vis_r5_o[25] : Qjc775);
assign Kyu675 = (W9b775 ? vis_r4_o[25] : Qjc775);
assign Dyu675 = (G8b775 ? vis_r11_o[25] : Qjc775);
assign Wxu675 = (Z7b775 ? vis_r10_o[25] : Qjc775);
assign Pxu675 = (S7b775 ? vis_r9_o[25] : Qjc775);
assign Ixu675 = (L7b775 ? vis_r8_o[25] : Qjc775);
assign Bxu675 = (E7b775 ? vis_r3_o[25] : Qjc775);
assign Uwu675 = (X6b775 ? vis_r2_o[25] : Qjc775);
assign Nwu675 = (Gi1775 ? vis_r1_o[25] : Qjc775);
assign Gwu675 = (Sp0775 ? vis_r0_o[25] : Qjc775);
assign Qjc775 = (~(Xjc775 & Ekc775));
assign Ekc775 = (Lkc775 & Skc775);
assign Skc775 = (~(Gec775 | Tz1l85[25]));
assign Lkc775 = (~(Zkc775 | Glc775));
assign Zkc775 = (Nlc775 & Ity675);
assign Nlc775 = (Tr1l85 & Ifc775);
assign Xjc775 = (Ulc775 & Bmc775);
assign Ulc775 = (Imc775 & Pmc775);
assign Pmc775 = (Cdb775 | Wmc775);
assign Imc775 = (~(Mbb775 & Sy1l85[25]));
assign Zvu675 = (Szb775 ? Dnc775 : vis_psp_o[22]);
assign Svu675 = (Zzb775 ? Dnc775 : vis_msp_o[22]);
assign Lvu675 = (N8b775 ? vis_r14_o[24] : Dnc775);
assign Evu675 = (U8b775 ? vis_r12_o[24] : Dnc775);
assign Xuu675 = (B9b775 ? vis_r7_o[24] : Dnc775);
assign Quu675 = (I9b775 ? vis_r6_o[24] : Dnc775);
assign Juu675 = (P9b775 ? vis_r5_o[24] : Dnc775);
assign Cuu675 = (W9b775 ? vis_r4_o[24] : Dnc775);
assign Vtu675 = (G8b775 ? vis_r11_o[24] : Dnc775);
assign Otu675 = (Z7b775 ? vis_r10_o[24] : Dnc775);
assign Htu675 = (S7b775 ? vis_r9_o[24] : Dnc775);
assign Atu675 = (L7b775 ? vis_r8_o[24] : Dnc775);
assign Tsu675 = (E7b775 ? vis_r3_o[24] : Dnc775);
assign Msu675 = (X6b775 ? vis_r2_o[24] : Dnc775);
assign Fsu675 = (Gi1775 ? vis_r1_o[24] : Dnc775);
assign Yru675 = (Sp0775 ? vis_r0_o[24] : Dnc775);
assign Dnc775 = (~(O90775 & Knc775));
assign Rru675 = (~(Rnc775 & Ync775));
assign Ync775 = (Foc775 | H20775);
assign Rnc775 = (Moc775 & Toc775);
assign Toc775 = (~(vis_pc_o[5] & Y00775));
assign Moc775 = (~(T10775 & haddr_o[6]));
assign Kru675 = (Szb775 ? Apc775 : vis_psp_o[4]);
assign Dru675 = (Zzb775 ? Apc775 : vis_msp_o[4]);
assign Wqu675 = (N8b775 ? vis_r14_o[6] : Apc775);
assign Pqu675 = (U8b775 ? vis_r12_o[6] : Apc775);
assign Iqu675 = (B9b775 ? vis_r7_o[6] : Apc775);
assign Bqu675 = (I9b775 ? vis_r6_o[6] : Apc775);
assign Upu675 = (P9b775 ? vis_r5_o[6] : Apc775);
assign Npu675 = (W9b775 ? vis_r4_o[6] : Apc775);
assign Gpu675 = (G8b775 ? vis_r11_o[6] : Apc775);
assign Zou675 = (Z7b775 ? vis_r10_o[6] : Apc775);
assign Sou675 = (S7b775 ? vis_r9_o[6] : Apc775);
assign Lou675 = (L7b775 ? vis_r8_o[6] : Apc775);
assign Eou675 = (E7b775 ? vis_r3_o[6] : Apc775);
assign Xnu675 = (X6b775 ? vis_r2_o[6] : Apc775);
assign Qnu675 = (Gi1775 ? vis_r1_o[6] : Apc775);
assign Jnu675 = (Sp0775 ? vis_r0_o[6] : Apc775);
assign Apc775 = (~(Hpc775 & Opc775));
assign Opc775 = (Vpc775 & Cqc775);
assign Cqc775 = (~(Gec775 | Tz1l85[6]));
assign Vpc775 = (~(Jqc775 | Qqc775));
assign Jqc775 = (Xqc775 & Apy675);
assign Xqc775 = (Dq1l85 & Ifc775);
assign Hpc775 = (Erc775 & Lrc775);
assign Erc775 = (Src775 & Zrc775);
assign Zrc775 = (Cdb775 | Gsc775);
assign Src775 = (~(Mbb775 & Sy1l85[6]));
assign Cnu675 = (~(Nsc775 & Usc775));
assign Usc775 = (Btc775 & Itc775);
assign Itc775 = (~(R00775 & vis_ipsr_o[5]));
assign Btc775 = (~(vis_pc_o[4] & Y00775));
assign Nsc775 = (Ptc775 & Wtc775);
assign Wtc775 = (~(T10775 & haddr_o[5]));
assign Ptc775 = (Duc775 | H20775);
assign Vmu675 = (Szb775 ? Kuc775 : vis_psp_o[3]);
assign Omu675 = (Zzb775 ? Kuc775 : vis_msp_o[3]);
assign Hmu675 = (N8b775 ? vis_r14_o[5] : Kuc775);
assign Amu675 = (U8b775 ? vis_r12_o[5] : Kuc775);
assign Tlu675 = (B9b775 ? vis_r7_o[5] : Kuc775);
assign Mlu675 = (I9b775 ? vis_r6_o[5] : Kuc775);
assign Flu675 = (P9b775 ? vis_r5_o[5] : Kuc775);
assign Yku675 = (W9b775 ? vis_r4_o[5] : Kuc775);
assign Rku675 = (G8b775 ? vis_r11_o[5] : Kuc775);
assign Kku675 = (Z7b775 ? vis_r10_o[5] : Kuc775);
assign Dku675 = (S7b775 ? vis_r9_o[5] : Kuc775);
assign Wju675 = (L7b775 ? vis_r8_o[5] : Kuc775);
assign Pju675 = (E7b775 ? vis_r3_o[5] : Kuc775);
assign Iju675 = (X6b775 ? vis_r2_o[5] : Kuc775);
assign Bju675 = (Gi1775 ? vis_r1_o[5] : Kuc775);
assign Uiu675 = (Sp0775 ? vis_r0_o[5] : Kuc775);
assign Kuc775 = (~(Mv5775 & Ruc775));
assign Niu675 = (~(Yuc775 & Fvc775));
assign Fvc775 = (Mvc775 & Tvc775);
assign Tvc775 = (~(R00775 & vis_ipsr_o[4]));
assign Mvc775 = (~(vis_pc_o[3] & Y00775));
assign Yuc775 = (Awc775 & Hwc775);
assign Hwc775 = (Jkb775 | Avz675);
assign Avz675 = (!haddr_o[4]);
assign Awc775 = (Owc775 | H20775);
assign Giu675 = (Szb775 ? Vwc775 : vis_psp_o[2]);
assign Zhu675 = (Zzb775 ? Vwc775 : vis_msp_o[2]);
assign Shu675 = (N8b775 ? vis_r14_o[4] : Vwc775);
assign Lhu675 = (U8b775 ? vis_r12_o[4] : Vwc775);
assign Ehu675 = (B9b775 ? vis_r7_o[4] : Vwc775);
assign Xgu675 = (I9b775 ? vis_r6_o[4] : Vwc775);
assign Qgu675 = (P9b775 ? vis_r5_o[4] : Vwc775);
assign Jgu675 = (W9b775 ? vis_r4_o[4] : Vwc775);
assign Cgu675 = (G8b775 ? vis_r11_o[4] : Vwc775);
assign Vfu675 = (Z7b775 ? vis_r10_o[4] : Vwc775);
assign Ofu675 = (S7b775 ? vis_r9_o[4] : Vwc775);
assign Hfu675 = (L7b775 ? vis_r8_o[4] : Vwc775);
assign Afu675 = (E7b775 ? vis_r3_o[4] : Vwc775);
assign Teu675 = (X6b775 ? vis_r2_o[4] : Vwc775);
assign Meu675 = (Gi1775 ? vis_r1_o[4] : Vwc775);
assign Feu675 = (Sp0775 ? vis_r0_o[4] : Vwc775);
assign Vwc775 = (~(Oh6775 & Cxc775));
assign Ydu675 = (~(Jxc775 & Qxc775));
assign Qxc775 = (Xxc775 & Eyc775);
assign Eyc775 = (Jkb775 | Isz675);
assign Isz675 = (!haddr_o[3]);
assign haddr_o[3] = (~(Lyc775 & Syc775));
assign Syc775 = (Jjc775 | Vpy675);
assign Lyc775 = (Zyc775 & Gzc775);
assign Gzc775 = (~(Nx1l85[2] & Dp3775));
assign Zyc775 = (~(Sy1l85[3] & Ms8775));
assign Xxc775 = (~(R00775 & vis_ipsr_o[3]));
assign Jxc775 = (Nzc775 & Uzc775);
assign Uzc775 = (~(Y00775 & vis_pc_o[2]));
assign Nzc775 = (~(Gpl675 & Ht8775));
assign Rdu675 = (Szb775 ? B0d775 : vis_psp_o[1]);
assign Kdu675 = (Zzb775 ? B0d775 : vis_msp_o[1]);
assign Ddu675 = (N8b775 ? vis_r14_o[3] : B0d775);
assign Wcu675 = (U8b775 ? vis_r12_o[3] : B0d775);
assign Pcu675 = (B9b775 ? vis_r7_o[3] : B0d775);
assign Icu675 = (I9b775 ? vis_r6_o[3] : B0d775);
assign Bcu675 = (P9b775 ? vis_r5_o[3] : B0d775);
assign Ubu675 = (W9b775 ? vis_r4_o[3] : B0d775);
assign Nbu675 = (G8b775 ? vis_r11_o[3] : B0d775);
assign Gbu675 = (Z7b775 ? vis_r10_o[3] : B0d775);
assign Zau675 = (S7b775 ? vis_r9_o[3] : B0d775);
assign Sau675 = (L7b775 ? vis_r8_o[3] : B0d775);
assign Lau675 = (E7b775 ? vis_r3_o[3] : B0d775);
assign Eau675 = (X6b775 ? vis_r2_o[3] : B0d775);
assign X9u675 = (Gi1775 ? vis_r1_o[3] : B0d775);
assign Q9u675 = (Sp0775 ? vis_r0_o[3] : B0d775);
assign B0d775 = (~(I0d775 & P0d775));
assign P0d775 = (W0d775 & D1d775);
assign D1d775 = (Cdb775 | K1d775);
assign W0d775 = (R1d775 & Y1d775);
assign Y1d775 = (~(F2d775 & F2s675));
assign F2d775 = (~(Ocb775 | M2d775));
assign R1d775 = (M3c775 | Pnb775);
assign I0d775 = (T2d775 & Sx6775);
assign T2d775 = (A3d775 & H3d775);
assign H3d775 = (~(Mbb775 & Sy1l85[3]));
assign J9u675 = (U41775 ? O3d775 : M62l85[1]);
assign U41775 = (!Mq3775);
assign Mq3775 = (~(hready_i & hprot_o[0]));
assign C9u675 = (~(V3d775 & C4d775));
assign C4d775 = (J4d775 | H20775);
assign V3d775 = (Q4d775 & X4d775);
assign X4d775 = (~(vis_pc_o[21] & Y00775));
assign Q4d775 = (~(T10775 & haddr_o[22]));
assign V8u675 = (Szb775 ? E5d775 : vis_psp_o[20]);
assign O8u675 = (Zzb775 ? E5d775 : vis_msp_o[20]);
assign H8u675 = (N8b775 ? vis_r14_o[22] : E5d775);
assign A8u675 = (U8b775 ? vis_r12_o[22] : E5d775);
assign T7u675 = (B9b775 ? vis_r7_o[22] : E5d775);
assign M7u675 = (I9b775 ? vis_r6_o[22] : E5d775);
assign F7u675 = (P9b775 ? vis_r5_o[22] : E5d775);
assign Y6u675 = (W9b775 ? vis_r4_o[22] : E5d775);
assign R6u675 = (G8b775 ? vis_r11_o[22] : E5d775);
assign K6u675 = (Z7b775 ? vis_r10_o[22] : E5d775);
assign D6u675 = (S7b775 ? vis_r9_o[22] : E5d775);
assign W5u675 = (L7b775 ? vis_r8_o[22] : E5d775);
assign P5u675 = (E7b775 ? vis_r3_o[22] : E5d775);
assign I5u675 = (X6b775 ? vis_r2_o[22] : E5d775);
assign B5u675 = (Gi1775 ? vis_r1_o[22] : E5d775);
assign U4u675 = (Sp0775 ? vis_r0_o[22] : E5d775);
assign E5d775 = (~(L5d775 & S5d775));
assign S5d775 = (Z5d775 & G6d775);
assign G6d775 = (~(N6d775 | Tz1l85[22]));
assign Z5d775 = (U6d775 & B7d775);
assign B7d775 = (~(I7d775 & Duy675));
assign I7d775 = (Uv1l85 & Ifc775);
assign U6d775 = (Cdb775 | P7d775);
assign L5d775 = (W7d775 & D8d775);
assign W7d775 = (K8d775 & R8d775);
assign R8d775 = (~(Mbb775 & Sy1l85[22]));
assign N4u675 = (~(Y8d775 & F9d775));
assign F9d775 = (M9d775 | H20775);
assign Y8d775 = (T9d775 & Aad775);
assign Aad775 = (~(vis_pc_o[20] & Y00775));
assign T9d775 = (~(T10775 & haddr_o[21]));
assign G4u675 = (Szb775 ? Had775 : vis_psp_o[19]);
assign Z3u675 = (Zzb775 ? Had775 : vis_msp_o[19]);
assign S3u675 = (N8b775 ? vis_r14_o[21] : Had775);
assign L3u675 = (U8b775 ? vis_r12_o[21] : Had775);
assign E3u675 = (B9b775 ? vis_r7_o[21] : Had775);
assign X2u675 = (I9b775 ? vis_r6_o[21] : Had775);
assign Q2u675 = (P9b775 ? vis_r5_o[21] : Had775);
assign J2u675 = (W9b775 ? vis_r4_o[21] : Had775);
assign C2u675 = (G8b775 ? vis_r11_o[21] : Had775);
assign V1u675 = (Z7b775 ? vis_r10_o[21] : Had775);
assign O1u675 = (S7b775 ? vis_r9_o[21] : Had775);
assign H1u675 = (L7b775 ? vis_r8_o[21] : Had775);
assign A1u675 = (E7b775 ? vis_r3_o[21] : Had775);
assign T0u675 = (X6b775 ? vis_r2_o[21] : Had775);
assign M0u675 = (Gi1775 ? vis_r1_o[21] : Had775);
assign F0u675 = (Sp0775 ? vis_r0_o[21] : Had775);
assign Had775 = (~(Oad775 & Vad775));
assign Vad775 = (Cbd775 & Jbd775);
assign Jbd775 = (~(Qbd775 | Tz1l85[21]));
assign Cbd775 = (Xbd775 & Ecd775);
assign Ecd775 = (~(Lcd775 & Kuy675));
assign Lcd775 = (Nv1l85 & Ifc775);
assign Xbd775 = (Cdb775 | Scd775);
assign Oad775 = (Zcd775 & Gdd775);
assign Zcd775 = (K8d775 & Ndd775);
assign Ndd775 = (~(Mbb775 & Sy1l85[21]));
assign Yzt675 = (~(Udd775 & Bed775));
assign Bed775 = (Ied775 | H20775);
assign Udd775 = (Ped775 & Wed775);
assign Wed775 = (~(vis_pc_o[19] & Y00775));
assign Ped775 = (~(T10775 & haddr_o[20]));
assign Rzt675 = (Szb775 ? Dfd775 : vis_psp_o[18]);
assign Kzt675 = (Zzb775 ? Dfd775 : vis_msp_o[18]);
assign Dzt675 = (N8b775 ? vis_r14_o[20] : Dfd775);
assign Wyt675 = (U8b775 ? vis_r12_o[20] : Dfd775);
assign Pyt675 = (B9b775 ? vis_r7_o[20] : Dfd775);
assign Iyt675 = (I9b775 ? vis_r6_o[20] : Dfd775);
assign Byt675 = (P9b775 ? vis_r5_o[20] : Dfd775);
assign Uxt675 = (W9b775 ? vis_r4_o[20] : Dfd775);
assign Nxt675 = (G8b775 ? vis_r11_o[20] : Dfd775);
assign Gxt675 = (Z7b775 ? vis_r10_o[20] : Dfd775);
assign Zwt675 = (S7b775 ? vis_r9_o[20] : Dfd775);
assign Swt675 = (L7b775 ? vis_r8_o[20] : Dfd775);
assign Lwt675 = (E7b775 ? vis_r3_o[20] : Dfd775);
assign Ewt675 = (X6b775 ? vis_r2_o[20] : Dfd775);
assign Xvt675 = (Gi1775 ? vis_r1_o[20] : Dfd775);
assign Qvt675 = (Sp0775 ? vis_r0_o[20] : Dfd775);
assign Dfd775 = (~(Kfd775 & Rfd775));
assign Rfd775 = (Yfd775 & Fgd775);
assign Fgd775 = (~(Mgd775 | Tz1l85[20]));
assign Yfd775 = (Tgd775 & Ahd775);
assign Ahd775 = (~(Hhd775 & Ruy675));
assign Hhd775 = (Bw1l85 & Ifc775);
assign Tgd775 = (Cdb775 | Ohd775);
assign Kfd775 = (Vhd775 & Cid775);
assign Vhd775 = (K8d775 & Jid775);
assign Jid775 = (~(Mbb775 & Sy1l85[20]));
assign Jvt675 = (~(Qid775 & Xid775));
assign Xid775 = (Ejd775 | H20775);
assign Qid775 = (Ljd775 & Sjd775);
assign Sjd775 = (~(vis_pc_o[18] & Y00775));
assign Ljd775 = (~(T10775 & haddr_o[19]));
assign Cvt675 = (Szb775 ? Zjd775 : vis_psp_o[17]);
assign Vut675 = (Zzb775 ? Zjd775 : vis_msp_o[17]);
assign Out675 = (N8b775 ? vis_r14_o[19] : Zjd775);
assign Hut675 = (U8b775 ? vis_r12_o[19] : Zjd775);
assign Aut675 = (B9b775 ? vis_r7_o[19] : Zjd775);
assign Ttt675 = (I9b775 ? vis_r6_o[19] : Zjd775);
assign Mtt675 = (P9b775 ? vis_r5_o[19] : Zjd775);
assign Ftt675 = (W9b775 ? vis_r4_o[19] : Zjd775);
assign Yst675 = (G8b775 ? vis_r11_o[19] : Zjd775);
assign Rst675 = (Z7b775 ? vis_r10_o[19] : Zjd775);
assign Kst675 = (S7b775 ? vis_r9_o[19] : Zjd775);
assign Dst675 = (L7b775 ? vis_r8_o[19] : Zjd775);
assign Wrt675 = (E7b775 ? vis_r3_o[19] : Zjd775);
assign Prt675 = (X6b775 ? vis_r2_o[19] : Zjd775);
assign Irt675 = (Gi1775 ? vis_r1_o[19] : Zjd775);
assign Brt675 = (Sp0775 ? vis_r0_o[19] : Zjd775);
assign Zjd775 = (~(Gkd775 & Nkd775));
assign Nkd775 = (Ukd775 & Bld775);
assign Bld775 = (~(Ild775 | Tz1l85[19]));
assign Ukd775 = (Pld775 & Wld775);
assign Wld775 = (~(Dmd775 & Fvy675));
assign Dmd775 = (Gv1l85 & Ifc775);
assign Pld775 = (Cdb775 | Kmd775);
assign Gkd775 = (Rmd775 & Ymd775);
assign Rmd775 = (K8d775 & Fnd775);
assign Fnd775 = (~(Mbb775 & Sy1l85[19]));
assign Uqt675 = (~(Mnd775 & Tnd775));
assign Tnd775 = (Aod775 | H20775);
assign Mnd775 = (Hod775 & Ood775);
assign Ood775 = (~(vis_pc_o[17] & Y00775));
assign Hod775 = (~(T10775 & haddr_o[18]));
assign Nqt675 = (Szb775 ? Vod775 : vis_psp_o[16]);
assign Gqt675 = (Zzb775 ? Vod775 : vis_msp_o[16]);
assign Zpt675 = (N8b775 ? vis_r14_o[18] : Vod775);
assign Spt675 = (U8b775 ? vis_r12_o[18] : Vod775);
assign Lpt675 = (B9b775 ? vis_r7_o[18] : Vod775);
assign Ept675 = (I9b775 ? vis_r6_o[18] : Vod775);
assign Xot675 = (P9b775 ? vis_r5_o[18] : Vod775);
assign Qot675 = (W9b775 ? vis_r4_o[18] : Vod775);
assign Jot675 = (G8b775 ? vis_r11_o[18] : Vod775);
assign Cot675 = (Z7b775 ? vis_r10_o[18] : Vod775);
assign Vnt675 = (S7b775 ? vis_r9_o[18] : Vod775);
assign Ont675 = (L7b775 ? vis_r8_o[18] : Vod775);
assign Hnt675 = (E7b775 ? vis_r3_o[18] : Vod775);
assign Ant675 = (X6b775 ? vis_r2_o[18] : Vod775);
assign Tmt675 = (Gi1775 ? vis_r1_o[18] : Vod775);
assign Mmt675 = (Sp0775 ? vis_r0_o[18] : Vod775);
assign Vod775 = (~(Cpd775 & Jpd775));
assign Jpd775 = (Qpd775 & Xpd775);
assign Xpd775 = (~(Eqd775 | Tz1l85[18]));
assign Qpd775 = (Lqd775 & Sqd775);
assign Sqd775 = (~(Zqd775 & Mvy675));
assign Zqd775 = (Zu1l85 & Ifc775);
assign Lqd775 = (Cdb775 | Grd775);
assign Cpd775 = (Nrd775 & Urd775);
assign Nrd775 = (K8d775 & Bsd775);
assign Bsd775 = (~(Mbb775 & Sy1l85[18]));
assign Fmt675 = (~(Isd775 & Psd775));
assign Psd775 = (Wsd775 | H20775);
assign Isd775 = (Dtd775 & Ktd775);
assign Ktd775 = (~(vis_pc_o[16] & Y00775));
assign Dtd775 = (~(T10775 & haddr_o[17]));
assign Ylt675 = (Szb775 ? Rtd775 : vis_psp_o[15]);
assign Rlt675 = (Zzb775 ? Rtd775 : vis_msp_o[15]);
assign Klt675 = (N8b775 ? vis_r14_o[17] : Rtd775);
assign Dlt675 = (U8b775 ? vis_r12_o[17] : Rtd775);
assign Wkt675 = (B9b775 ? vis_r7_o[17] : Rtd775);
assign Pkt675 = (I9b775 ? vis_r6_o[17] : Rtd775);
assign Ikt675 = (P9b775 ? vis_r5_o[17] : Rtd775);
assign Bkt675 = (W9b775 ? vis_r4_o[17] : Rtd775);
assign Ujt675 = (G8b775 ? vis_r11_o[17] : Rtd775);
assign Njt675 = (Z7b775 ? vis_r10_o[17] : Rtd775);
assign Gjt675 = (S7b775 ? vis_r9_o[17] : Rtd775);
assign Zit675 = (L7b775 ? vis_r8_o[17] : Rtd775);
assign Sit675 = (E7b775 ? vis_r3_o[17] : Rtd775);
assign Lit675 = (X6b775 ? vis_r2_o[17] : Rtd775);
assign Eit675 = (Gi1775 ? vis_r1_o[17] : Rtd775);
assign Xht675 = (Sp0775 ? vis_r0_o[17] : Rtd775);
assign Rtd775 = (~(Ytd775 & Fud775));
assign Fud775 = (Mud775 & Tud775);
assign Tud775 = (Avd775 & Hvd775);
assign Mud775 = (Ovd775 & Vvd775);
assign Vvd775 = (~(Cwd775 & Tvy675));
assign Cwd775 = (Lu1l85 & Ifc775);
assign Ovd775 = (Cdb775 | Jwd775);
assign Ytd775 = (Qwd775 & Xwd775);
assign Qwd775 = (K8d775 & Exd775);
assign Exd775 = (~(Mbb775 & Sy1l85[17]));
assign Qht675 = (~(Lxd775 & Sxd775));
assign Sxd775 = (Zxd775 | H20775);
assign Lxd775 = (Gyd775 & Nyd775);
assign Nyd775 = (~(vis_pc_o[15] & Y00775));
assign Gyd775 = (~(T10775 & haddr_o[16]));
assign haddr_o[16] = (~(Uyd775 & Bzd775));
assign Bzd775 = (~(Nx1l85[15] & Dp3775));
assign Uyd775 = (Izd775 & Pzd775);
assign Pzd775 = (Jjc775 | Awy675);
assign Izd775 = (~(Sy1l85[16] & Ms8775));
assign Jht675 = (Szb775 ? Wzd775 : vis_psp_o[14]);
assign Cht675 = (Zzb775 ? Wzd775 : vis_msp_o[14]);
assign Vgt675 = (N8b775 ? vis_r14_o[16] : Wzd775);
assign Ogt675 = (U8b775 ? vis_r12_o[16] : Wzd775);
assign Hgt675 = (B9b775 ? vis_r7_o[16] : Wzd775);
assign Agt675 = (I9b775 ? vis_r6_o[16] : Wzd775);
assign Tft675 = (P9b775 ? vis_r5_o[16] : Wzd775);
assign Mft675 = (W9b775 ? vis_r4_o[16] : Wzd775);
assign Fft675 = (G8b775 ? vis_r11_o[16] : Wzd775);
assign Yet675 = (Z7b775 ? vis_r10_o[16] : Wzd775);
assign Ret675 = (S7b775 ? vis_r9_o[16] : Wzd775);
assign Ket675 = (L7b775 ? vis_r8_o[16] : Wzd775);
assign Det675 = (E7b775 ? vis_r3_o[16] : Wzd775);
assign Wdt675 = (X6b775 ? vis_r2_o[16] : Wzd775);
assign Pdt675 = (Gi1775 ? vis_r1_o[16] : Wzd775);
assign Idt675 = (Sp0775 ? vis_r0_o[16] : Wzd775);
assign Wzd775 = (~(D0e775 & K0e775));
assign K0e775 = (R0e775 & Y0e775);
assign Y0e775 = (~(F1e775 | Tz1l85[16]));
assign R0e775 = (M1e775 & T1e775);
assign T1e775 = (~(A2e775 & Awy675));
assign A2e775 = (Eu1l85 & Ifc775);
assign M1e775 = (Cdb775 | H2e775);
assign D0e775 = (O2e775 & V2e775);
assign O2e775 = (K8d775 & C3e775);
assign C3e775 = (~(Mbb775 & Sy1l85[16]));
assign K8d775 = (J3e775 & M3c775);
assign Bdt675 = (~(Q3e775 & X3e775));
assign X3e775 = (E4e775 | H20775);
assign Q3e775 = (L4e775 & S4e775);
assign S4e775 = (~(vis_pc_o[13] & Y00775));
assign L4e775 = (~(T10775 & haddr_o[14]));
assign Uct675 = (Szb775 ? Z4e775 : vis_psp_o[12]);
assign Nct675 = (Zzb775 ? Z4e775 : vis_msp_o[12]);
assign Gct675 = (N8b775 ? vis_r14_o[14] : Z4e775);
assign Zbt675 = (U8b775 ? vis_r12_o[14] : Z4e775);
assign Sbt675 = (B9b775 ? vis_r7_o[14] : Z4e775);
assign Lbt675 = (I9b775 ? vis_r6_o[14] : Z4e775);
assign Ebt675 = (P9b775 ? vis_r5_o[14] : Z4e775);
assign Xat675 = (W9b775 ? vis_r4_o[14] : Z4e775);
assign Qat675 = (G8b775 ? vis_r11_o[14] : Z4e775);
assign Jat675 = (Z7b775 ? vis_r10_o[14] : Z4e775);
assign Cat675 = (S7b775 ? vis_r9_o[14] : Z4e775);
assign V9t675 = (L7b775 ? vis_r8_o[14] : Z4e775);
assign O9t675 = (E7b775 ? vis_r3_o[14] : Z4e775);
assign H9t675 = (X6b775 ? vis_r2_o[14] : Z4e775);
assign A9t675 = (Gi1775 ? vis_r1_o[14] : Z4e775);
assign T8t675 = (Sp0775 ? vis_r0_o[14] : Z4e775);
assign Z4e775 = (~(G5e775 & N5e775));
assign N5e775 = (U5e775 & B6e775);
assign B6e775 = (~(I6e775 | Tz1l85[14]));
assign U5e775 = (P6e775 & W6e775);
assign W6e775 = (~(D7e775 & Owy675));
assign D7e775 = (Xt1l85 & Ifc775);
assign P6e775 = (Cdb775 | K7e775);
assign G5e775 = (R7e775 & Y7e775);
assign R7e775 = (F8e775 & M8e775);
assign M8e775 = (~(Mbb775 & Sy1l85[14]));
assign M8t675 = (~(T8e775 & A9e775));
assign A9e775 = (H9e775 | H20775);
assign T8e775 = (O9e775 & V9e775);
assign V9e775 = (~(vis_pc_o[12] & Y00775));
assign O9e775 = (~(T10775 & haddr_o[13]));
assign F8t675 = (Szb775 ? Cae775 : vis_psp_o[11]);
assign Y7t675 = (Zzb775 ? Cae775 : vis_msp_o[11]);
assign R7t675 = (N8b775 ? vis_r14_o[13] : Cae775);
assign K7t675 = (U8b775 ? vis_r12_o[13] : Cae775);
assign D7t675 = (B9b775 ? vis_r7_o[13] : Cae775);
assign W6t675 = (I9b775 ? vis_r6_o[13] : Cae775);
assign P6t675 = (P9b775 ? vis_r5_o[13] : Cae775);
assign I6t675 = (W9b775 ? vis_r4_o[13] : Cae775);
assign B6t675 = (G8b775 ? vis_r11_o[13] : Cae775);
assign U5t675 = (Z7b775 ? vis_r10_o[13] : Cae775);
assign N5t675 = (S7b775 ? vis_r9_o[13] : Cae775);
assign G5t675 = (L7b775 ? vis_r8_o[13] : Cae775);
assign Z4t675 = (E7b775 ? vis_r3_o[13] : Cae775);
assign S4t675 = (X6b775 ? vis_r2_o[13] : Cae775);
assign L4t675 = (Gi1775 ? vis_r1_o[13] : Cae775);
assign E4t675 = (Sp0775 ? vis_r0_o[13] : Cae775);
assign Cae775 = (~(Jae775 & Qae775));
assign Qae775 = (Xae775 & Ebe775);
assign Ebe775 = (~(Lbe775 | Tz1l85[13]));
assign Xae775 = (Sbe775 & Zbe775);
assign Zbe775 = (~(Gce775 & Vwy675));
assign Gce775 = (Qt1l85 & Ifc775);
assign Sbe775 = (Cdb775 | Nce775);
assign Jae775 = (Uce775 & Bde775);
assign Uce775 = (F8e775 & Ide775);
assign Ide775 = (~(Mbb775 & Sy1l85[13]));
assign X3t675 = (~(Pde775 & Wde775));
assign Wde775 = (Dee775 | H20775);
assign Pde775 = (Kee775 & Ree775);
assign Ree775 = (~(vis_pc_o[11] & Y00775));
assign Kee775 = (~(T10775 & haddr_o[12]));
assign haddr_o[12] = (~(Yee775 & Ffe775));
assign Ffe775 = (~(Nx1l85[11] & Dp3775));
assign Yee775 = (Mfe775 & Tfe775);
assign Tfe775 = (Jjc775 | Cxy675);
assign Mfe775 = (~(Sy1l85[12] & Ms8775));
assign Q3t675 = (Szb775 ? Age775 : vis_psp_o[10]);
assign J3t675 = (Zzb775 ? Age775 : vis_msp_o[10]);
assign C3t675 = (N8b775 ? vis_r14_o[12] : Age775);
assign V2t675 = (U8b775 ? vis_r12_o[12] : Age775);
assign O2t675 = (B9b775 ? vis_r7_o[12] : Age775);
assign H2t675 = (I9b775 ? vis_r6_o[12] : Age775);
assign A2t675 = (P9b775 ? vis_r5_o[12] : Age775);
assign T1t675 = (W9b775 ? vis_r4_o[12] : Age775);
assign M1t675 = (G8b775 ? vis_r11_o[12] : Age775);
assign F1t675 = (Z7b775 ? vis_r10_o[12] : Age775);
assign Y0t675 = (S7b775 ? vis_r9_o[12] : Age775);
assign R0t675 = (L7b775 ? vis_r8_o[12] : Age775);
assign K0t675 = (E7b775 ? vis_r3_o[12] : Age775);
assign D0t675 = (X6b775 ? vis_r2_o[12] : Age775);
assign Wzs675 = (Gi1775 ? vis_r1_o[12] : Age775);
assign Pzs675 = (Sp0775 ? vis_r0_o[12] : Age775);
assign Age775 = (~(Hge775 & Oge775));
assign Oge775 = (Vge775 & Che775);
assign Che775 = (~(Jhe775 | Tz1l85[12]));
assign Vge775 = (Qhe775 & Xhe775);
assign Xhe775 = (~(Eie775 & Cxy675));
assign Eie775 = (Jt1l85 & Ifc775);
assign Qhe775 = (Cdb775 | Lie775);
assign Hge775 = (Sie775 & Zie775);
assign Sie775 = (F8e775 & Gje775);
assign Gje775 = (~(Mbb775 & Sy1l85[12]));
assign Izs675 = (~(Nje775 & Uje775));
assign Uje775 = (Bke775 | H20775);
assign Nje775 = (Ike775 & Pke775);
assign Pke775 = (~(T10775 & haddr_o[11]));
assign haddr_o[11] = (~(Wke775 & Dle775));
assign Dle775 = (Jjc775 | Jxy675);
assign Wke775 = (Kle775 & Rle775);
assign Rle775 = (~(Nx1l85[10] & Dp3775));
assign Kle775 = (~(Sy1l85[11] & Ms8775));
assign Ike775 = (~(vis_pc_o[10] & Y00775));
assign Bzs675 = (Szb775 ? Yle775 : vis_psp_o[9]);
assign Uys675 = (Zzb775 ? Yle775 : vis_msp_o[9]);
assign Nys675 = (N8b775 ? vis_r14_o[11] : Yle775);
assign Gys675 = (U8b775 ? vis_r12_o[11] : Yle775);
assign Zxs675 = (B9b775 ? vis_r7_o[11] : Yle775);
assign Sxs675 = (I9b775 ? vis_r6_o[11] : Yle775);
assign Lxs675 = (P9b775 ? vis_r5_o[11] : Yle775);
assign Exs675 = (W9b775 ? vis_r4_o[11] : Yle775);
assign Xws675 = (G8b775 ? vis_r11_o[11] : Yle775);
assign Qws675 = (Z7b775 ? vis_r10_o[11] : Yle775);
assign Jws675 = (S7b775 ? vis_r9_o[11] : Yle775);
assign Cws675 = (L7b775 ? vis_r8_o[11] : Yle775);
assign Vvs675 = (E7b775 ? vis_r3_o[11] : Yle775);
assign Ovs675 = (X6b775 ? vis_r2_o[11] : Yle775);
assign Hvs675 = (Gi1775 ? vis_r1_o[11] : Yle775);
assign Avs675 = (Sp0775 ? vis_r0_o[11] : Yle775);
assign Yle775 = (~(Fme775 & Mme775));
assign Mme775 = (Tme775 & Ane775);
assign Ane775 = (Hne775 & One775);
assign Tme775 = (Vne775 & Coe775);
assign Coe775 = (~(Joe775 & Jxy675));
assign Joe775 = (~(Qoe775 | Ocb775));
assign Vne775 = (Cdb775 | Xoe775);
assign Fme775 = (Epe775 & Lpe775);
assign Epe775 = (F8e775 & Spe775);
assign Spe775 = (~(Mbb775 & Sy1l85[11]));
assign Tus675 = (~(Zpe775 & Gqe775));
assign Gqe775 = (Nqe775 | H20775);
assign Zpe775 = (Uqe775 & Bre775);
assign Bre775 = (~(vis_pc_o[9] & Y00775));
assign Uqe775 = (Jkb775 | Nkz675);
assign Nkz675 = (!haddr_o[10]);
assign Mus675 = (Szb775 ? Ire775 : vis_psp_o[8]);
assign Fus675 = (Zzb775 ? Ire775 : vis_msp_o[8]);
assign Yts675 = (N8b775 ? vis_r14_o[10] : Ire775);
assign Rts675 = (U8b775 ? vis_r12_o[10] : Ire775);
assign Kts675 = (B9b775 ? vis_r7_o[10] : Ire775);
assign Dts675 = (I9b775 ? vis_r6_o[10] : Ire775);
assign Wss675 = (P9b775 ? vis_r5_o[10] : Ire775);
assign Pss675 = (W9b775 ? vis_r4_o[10] : Ire775);
assign Iss675 = (G8b775 ? vis_r11_o[10] : Ire775);
assign Bss675 = (Z7b775 ? vis_r10_o[10] : Ire775);
assign Urs675 = (S7b775 ? vis_r9_o[10] : Ire775);
assign Nrs675 = (L7b775 ? vis_r8_o[10] : Ire775);
assign Grs675 = (E7b775 ? vis_r3_o[10] : Ire775);
assign Zqs675 = (X6b775 ? vis_r2_o[10] : Ire775);
assign Sqs675 = (Gi1775 ? vis_r1_o[10] : Ire775);
assign Lqs675 = (Sp0775 ? vis_r0_o[10] : Ire775);
assign Ire775 = (~(Pre775 & Wre775));
assign Pre775 = (Dse775 & Kse775);
assign Eqs675 = (Yse775 ? Rse775 : N6i675);
assign Yse775 = (Fte775 & hready_i);
assign Fte775 = (Zx6775 & Mte775);
assign Mte775 = (Tte775 | Sry675);
assign Rse775 = (Of8775 ? Xqy675 : Aue775);
assign Xps675 = (Szb775 ? Hue775 : vis_psp_o[0]);
assign Qps675 = (Zzb775 ? Hue775 : vis_msp_o[0]);
assign Jps675 = (N8b775 ? vis_r14_o[2] : Hue775);
assign Cps675 = (U8b775 ? vis_r12_o[2] : Hue775);
assign U8b775 = (!Oue775);
assign Vos675 = (B9b775 ? vis_r7_o[2] : Hue775);
assign B9b775 = (!Vue775);
assign Oos675 = (I9b775 ? vis_r6_o[2] : Hue775);
assign Hos675 = (P9b775 ? vis_r5_o[2] : Hue775);
assign P9b775 = (!Cve775);
assign Aos675 = (W9b775 ? vis_r4_o[2] : Hue775);
assign W9b775 = (!Jve775);
assign Tns675 = (G8b775 ? vis_r11_o[2] : Hue775);
assign G8b775 = (!Qve775);
assign Mns675 = (Z7b775 ? vis_r10_o[2] : Hue775);
assign Fns675 = (S7b775 ? vis_r9_o[2] : Hue775);
assign S7b775 = (!Xve775);
assign Yms675 = (L7b775 ? vis_r8_o[2] : Hue775);
assign L7b775 = (!Ewe775);
assign Rms675 = (E7b775 ? vis_r3_o[2] : Hue775);
assign E7b775 = (!Lwe775);
assign Kms675 = (X6b775 ? vis_r2_o[2] : Hue775);
assign Dms675 = (Gi1775 ? vis_r1_o[2] : Hue775);
assign Gi1775 = (!Swe775);
assign Wls675 = (Sp0775 ? vis_r0_o[2] : Hue775);
assign Sp0775 = (!Zwe775);
assign Hue775 = (~(T26775 & Gxe775));
assign Pls675 = (~(Nxe775 & Uxe775));
assign Uxe775 = (Bye775 & Iye775);
assign Iye775 = (~(T10775 & haddr_o[9]));
assign haddr_o[9] = (~(Pye775 & Wye775));
assign Wye775 = (Jjc775 | Yny675);
assign Pye775 = (Dze775 & Kze775);
assign Kze775 = (~(Nx1l85[8] & Dp3775));
assign Dze775 = (~(Sy1l85[9] & Ms8775));
assign Bye775 = (~(N6i675 & R00775));
assign Nxe775 = (Rze775 & Yze775);
assign Yze775 = (~(vis_pc_o[8] & Y00775));
assign Rze775 = (F0f775 | H20775);
assign Ils675 = (Szb775 ? M0f775 : vis_psp_o[7]);
assign Bls675 = (Zzb775 ? M0f775 : vis_msp_o[7]);
assign Uks675 = (N8b775 ? vis_r14_o[9] : M0f775);
assign Nks675 = (Oue775 ? M0f775 : vis_r12_o[9]);
assign Gks675 = (Vue775 ? M0f775 : vis_r7_o[9]);
assign Zjs675 = (I9b775 ? vis_r6_o[9] : M0f775);
assign Sjs675 = (Cve775 ? M0f775 : vis_r5_o[9]);
assign Ljs675 = (Jve775 ? M0f775 : vis_r4_o[9]);
assign Ejs675 = (Qve775 ? M0f775 : vis_r11_o[9]);
assign Xis675 = (Z7b775 ? vis_r10_o[9] : M0f775);
assign Qis675 = (Xve775 ? M0f775 : vis_r9_o[9]);
assign Jis675 = (Ewe775 ? M0f775 : vis_r8_o[9]);
assign Cis675 = (Lwe775 ? M0f775 : vis_r3_o[9]);
assign Vhs675 = (X6b775 ? vis_r2_o[9] : M0f775);
assign Ohs675 = (Swe775 ? M0f775 : vis_r1_o[9]);
assign Hhs675 = (Zwe775 ? M0f775 : vis_r0_o[9]);
assign M0f775 = (Aue775 | T0f775);
assign Ahs675 = (~(A1f775 & H1f775));
assign H1f775 = (O1f775 | H20775);
assign A1f775 = (V1f775 & C2f775);
assign C2f775 = (Jkb775 | I7z675);
assign I7z675 = (!haddr_o[8]);
assign haddr_o[8] = (~(J2f775 & Q2f775));
assign Q2f775 = (Jjc775 | Moy675);
assign J2f775 = (X2f775 & E3f775);
assign E3f775 = (~(Nx1l85[7] & Dp3775));
assign X2f775 = (~(Sy1l85[8] & Ms8775));
assign Jkb775 = (!T10775);
assign V1f775 = (~(vis_pc_o[7] & Y00775));
assign Tgs675 = (Szb775 ? L3f775 : vis_psp_o[6]);
assign Mgs675 = (Zzb775 ? L3f775 : vis_msp_o[6]);
assign Fgs675 = (N8b775 ? vis_r14_o[8] : L3f775);
assign Yfs675 = (Oue775 ? L3f775 : vis_r12_o[8]);
assign Rfs675 = (Vue775 ? L3f775 : vis_r7_o[8]);
assign Kfs675 = (I9b775 ? vis_r6_o[8] : L3f775);
assign Dfs675 = (Cve775 ? L3f775 : vis_r5_o[8]);
assign Wes675 = (Jve775 ? L3f775 : vis_r4_o[8]);
assign Pes675 = (Qve775 ? L3f775 : vis_r11_o[8]);
assign Ies675 = (Z7b775 ? vis_r10_o[8] : L3f775);
assign Bes675 = (Xve775 ? L3f775 : vis_r9_o[8]);
assign Uds675 = (Ewe775 ? L3f775 : vis_r8_o[8]);
assign Nds675 = (Lwe775 ? L3f775 : vis_r3_o[8]);
assign Gds675 = (X6b775 ? vis_r2_o[8] : L3f775);
assign Zcs675 = (Swe775 ? L3f775 : vis_r1_o[8]);
assign Scs675 = (Zwe775 ? L3f775 : vis_r0_o[8]);
assign L3f775 = (~(S3f775 & Z3f775));
assign Z3f775 = (G4f775 & N4f775);
assign N4f775 = (~(U4f775 | Tz1l85[8]));
assign G4f775 = (B5f775 & I5f775);
assign I5f775 = (~(P5f775 & Moy675));
assign P5f775 = (Wp1l85 & Ifc775);
assign B5f775 = (Cdb775 | W5f775);
assign S3f775 = (D6f775 & K6f775);
assign D6f775 = (F8e775 & R6f775);
assign R6f775 = (~(Mbb775 & Sy1l85[8]));
assign Lcs675 = (~(Y6f775 & F7f775));
assign F7f775 = (M7f775 | H20775);
assign Y6f775 = (T7f775 & A8f775);
assign A8f775 = (~(vis_pc_o[14] & Y00775));
assign T7f775 = (~(T10775 & haddr_o[15]));
assign Ecs675 = (Szb775 ? H8f775 : vis_psp_o[13]);
assign Xbs675 = (Zzb775 ? H8f775 : vis_msp_o[13]);
assign Qbs675 = (N8b775 ? vis_r14_o[15] : H8f775);
assign Jbs675 = (Oue775 ? H8f775 : vis_r12_o[15]);
assign Cbs675 = (Vue775 ? H8f775 : vis_r7_o[15]);
assign Vas675 = (I9b775 ? vis_r6_o[15] : H8f775);
assign Oas675 = (Cve775 ? H8f775 : vis_r5_o[15]);
assign Has675 = (Jve775 ? H8f775 : vis_r4_o[15]);
assign Aas675 = (Qve775 ? H8f775 : vis_r11_o[15]);
assign T9s675 = (Z7b775 ? vis_r10_o[15] : H8f775);
assign M9s675 = (Xve775 ? H8f775 : vis_r9_o[15]);
assign F9s675 = (Ewe775 ? H8f775 : vis_r8_o[15]);
assign Y8s675 = (Lwe775 ? H8f775 : vis_r3_o[15]);
assign R8s675 = (X6b775 ? vis_r2_o[15] : H8f775);
assign K8s675 = (Swe775 ? H8f775 : vis_r1_o[15]);
assign D8s675 = (Zwe775 ? H8f775 : vis_r0_o[15]);
assign H8f775 = (~(O8f775 & V8f775));
assign V8f775 = (C9f775 & J9f775);
assign J9f775 = (~(Q9f775 | Tz1l85[15]));
assign C9f775 = (X9f775 & Eaf775);
assign Eaf775 = (~(Laf775 & Hwy675));
assign Laf775 = (Su1l85 & Ifc775);
assign X9f775 = (Cdb775 | Saf775);
assign O8f775 = (Zaf775 & Gbf775);
assign Zaf775 = (F8e775 & Nbf775);
assign Nbf775 = (~(Mbb775 & Sy1l85[15]));
assign F8e775 = (~(Ubf775 | Gec775));
assign Ubf775 = (!Kse775);
assign W7s675 = (~(Bcf775 & Icf775));
assign Icf775 = (Pcf775 | H20775);
assign Bcf775 = (Wcf775 & Ddf775);
assign Ddf775 = (~(vis_pc_o[22] & Y00775));
assign Wcf775 = (~(T10775 & haddr_o[23]));
assign P7s675 = (Szb775 ? Kdf775 : vis_psp_o[21]);
assign Szb775 = (Rdf775 & Gum675);
assign Rdf775 = (!Ydf775);
assign I7s675 = (Zzb775 ? Kdf775 : vis_msp_o[21]);
assign Zzb775 = (~(Ydf775 | Gum675));
assign Ydf775 = (~(Fef775 & Mef775));
assign Fef775 = (Tef775 & Aff775);
assign B7s675 = (N8b775 ? vis_r14_o[23] : Kdf775);
assign N8b775 = (~(Hff775 & Off775));
assign U6s675 = (Oue775 ? Kdf775 : vis_r12_o[23]);
assign Oue775 = (Vff775 & Hff775);
assign Vff775 = (~(Cgf775 | Jgf775));
assign N6s675 = (Vue775 ? Kdf775 : vis_r7_o[23]);
assign Vue775 = (Qgf775 & Xgf775);
assign Qgf775 = (Tef775 & Ehf775);
assign G6s675 = (I9b775 ? vis_r6_o[23] : Kdf775);
assign I9b775 = (~(Hff775 & Xgf775));
assign Z5s675 = (Cve775 ? Kdf775 : vis_r5_o[23]);
assign Cve775 = (Lhf775 & Mef775);
assign Lhf775 = (Jgf775 & Tef775);
assign S5s675 = (Jve775 ? Kdf775 : vis_r4_o[23]);
assign Jve775 = (Shf775 & Hff775);
assign Hff775 = (Zhf775 & Tef775);
assign Shf775 = (~(Cgf775 | Aff775));
assign L5s675 = (Qve775 ? Kdf775 : vis_r11_o[23]);
assign Qve775 = (Gif775 & Off775);
assign E5s675 = (Z7b775 ? vis_r10_o[23] : Kdf775);
assign Z7b775 = (~(Off775 & Nif775));
assign Off775 = (~(Jgf775 | Uif775));
assign X4s675 = (Xve775 ? Kdf775 : vis_r9_o[23]);
assign Xve775 = (Bjf775 & Mef775);
assign Bjf775 = (~(Tef775 | Jgf775));
assign Q4s675 = (Ewe775 ? Kdf775 : vis_r8_o[23]);
assign Ewe775 = (Ijf775 & Uif775);
assign Ijf775 = (Nif775 & Aff775);
assign J4s675 = (Lwe775 ? Kdf775 : vis_r3_o[23]);
assign Lwe775 = (Gif775 & Xgf775);
assign Gif775 = (~(Tef775 | Zhf775));
assign C4s675 = (X6b775 ? vis_r2_o[23] : Kdf775);
assign X6b775 = (~(Xgf775 & Nif775));
assign Xgf775 = (~(Aff775 | Uif775));
assign V3s675 = (Swe775 ? Kdf775 : vis_r1_o[23]);
assign Swe775 = (Pjf775 & Mef775);
assign Mef775 = (~(Cgf775 | Zhf775));
assign Zhf775 = (!Ehf775);
assign Pjf775 = (~(Aff775 | Tef775));
assign O3s675 = (Zwe775 ? Kdf775 : vis_r0_o[23]);
assign Zwe775 = (Wjf775 & Uif775);
assign Uif775 = (!Cgf775);
assign Cgf775 = (Dkf775 | Kkf775);
assign Dkf775 = (~(hready_i & Rkf775));
assign Wjf775 = (Jgf775 & Nif775);
assign Nif775 = (~(Ehf775 | Tef775));
assign Tef775 = (~(Ykf775 & Flf775));
assign Flf775 = (Mlf775 & Tlf775);
assign Tlf775 = (Amf775 | Hmf775);
assign Mlf775 = (Omf775 & Vmf775);
assign Vmf775 = (Cnf775 | Jnf775);
assign Omf775 = (Qnf775 | Xnf775);
assign Ehf775 = (~(Eof775 & Lof775));
assign Lof775 = (Sof775 & Zof775);
assign Zof775 = (Gpf775 | Xnf775);
assign Sof775 = (Bx8775 | Hmf775);
assign Eof775 = (Npf775 & Upf775);
assign Upf775 = (Bqf775 | Jnf775);
assign Jgf775 = (!Aff775);
assign Aff775 = (~(Ykf775 & Iqf775));
assign Iqf775 = (Pqf775 & Wqf775);
assign Wqf775 = (Drf775 | Xnf775);
assign Pqf775 = (Krf775 & Rrf775);
assign Rrf775 = (Fd9775 | Hmf775);
assign Krf775 = (Yrf775 | Jnf775);
assign Ykf775 = (Npf775 & Fsf775);
assign Npf775 = (Msf775 & hready_i);
assign Msf775 = (Rkf775 & Tsf775);
assign Rkf775 = (~(Atf775 & Htf775));
assign Htf775 = (Otf775 & Vtf775);
assign Vtf775 = (Cuf775 & Juf775);
assign Juf775 = (~(Quf775 & Sh1775));
assign Quf775 = (~(Xuf775 | N0p675));
assign Cuf775 = (Evf775 & Lvf775);
assign Otf775 = (Svf775 & Zvf775);
assign Zvf775 = (~(Gwf775 & Nwf775));
assign Nwf775 = (Uwf775 | Bxf775);
assign Bxf775 = (Vxo675 ? Pxf775 : Ixf775);
assign Ixf775 = (~(Wxf775 & Dyf775));
assign Dyf775 = (Zry675 | Pw9775);
assign Uwf775 = (~(Kyf775 & Ryf775));
assign Kyf775 = (Yyf775 | D1z675);
assign Svf775 = (Fzf775 & Mzf775);
assign Mzf775 = (~(Mwo675 & Tzf775));
assign Tzf775 = (~(A0g775 & H0g775));
assign H0g775 = (~(O0g775 & V0g775));
assign A0g775 = (~(C1g775 & E5z675));
assign Fzf775 = (~(J1g775 & M71775));
assign J1g775 = (~(Q1g775 & X1g775));
assign X1g775 = (~(E2g775 & Dny675));
assign E2g775 = (~(L2g775 | X5p675));
assign Q1g775 = (S2g775 & Z2g775);
assign Z2g775 = (~(G3g775 & N3g775));
assign G3g775 = (~(U3g775 | Wxf775));
assign S2g775 = (~(B4g775 & Ub1775));
assign B4g775 = (N0p675 & Kny675);
assign Atf775 = (I4g775 & P4g775);
assign P4g775 = (W4g775 & D5g775);
assign D5g775 = (~(Os9775 & Nzy675));
assign W4g775 = (K5g775 & R5g775);
assign R5g775 = (~(Y5g775 & F6g775));
assign K5g775 = (~(V0g775 & M6g775));
assign I4g775 = (T6g775 & A7g775);
assign A7g775 = (F3p675 ? O7g775 : H7g775);
assign O7g775 = (~(V7g775 & Sfa775));
assign H7g775 = (C8g775 | Kp3775);
assign T6g775 = (J8g775 & Q8g775);
assign Q8g775 = (~(Qza775 & T5a775));
assign J8g775 = (Rto675 ? E9g775 : X8g775);
assign E9g775 = (L9g775 & S9g775);
assign S9g775 = (Yyf775 | C8g775);
assign L9g775 = (Z9g775 & Gag775);
assign Gag775 = (~(Nag775 & Uag775));
assign Nag775 = (~(Bbg775 | Ibg775));
assign Z9g775 = (~(F6g775 & Pbg775));
assign Pbg775 = (~(Wbg775 & Dcg775));
assign Dcg775 = (~(Kcg775 & Rcg775));
assign Kcg775 = (~(Vya775 | Zry675));
assign X8g775 = (Ycg775 & Fdg775);
assign Fdg775 = (~(Mdg775 & Tdg775));
assign Ycg775 = (Aeg775 & Heg775);
assign Heg775 = (~(Oeg775 & Uag775));
assign Oeg775 = (~(Veg775 | X5p675));
assign Aeg775 = (~(Cfg775 & M6g775));
assign Cfg775 = (Kny675 & Pw9775);
assign Kdf775 = (~(Jfg775 & Qfg775));
assign Jfg775 = (Xfg775 & J3e775);
assign H3s675 = (J5c775 ? Egg775 : vis_apsr_o[3]);
assign J5c775 = (hready_i & Lgg775);
assign Lgg775 = (~(Sgg775 & Br0775));
assign Egg775 = (~(Zgg775 & Ghg775));
assign Ghg775 = (D70775 | B1c775);
assign D70775 = (!Nhg775);
assign Zgg775 = (Uhg775 & Big775);
assign Big775 = (~(Br0775 & Iig775));
assign Br0775 = (~(Ys0775 | Nhg775));
assign Nhg775 = (Zx6775 & At1775);
assign Uhg775 = (~(Ys0775 & Pig775));
assign Ys0775 = (!Yz0775);
assign Yz0775 = (~(Wig775 & Inb775));
assign A3s675 = (~(Djg775 & Kjg775));
assign Kjg775 = (Rjg775 & Yjg775);
assign Yjg775 = (~(vis_apsr_o[3] & R00775));
assign R00775 = (~(Ht8775 | Lvf775));
assign Rjg775 = (~(Y00775 & vis_pc_o[30]));
assign Y00775 = (~(Ht8775 | Fkg775));
assign Djg775 = (Mkg775 & Tkg775);
assign Tkg775 = (~(T10775 & haddr_o[31]));
assign T10775 = (Alg775 & H20775);
assign Alg775 = (Hlg775 & Olg775);
assign Hlg775 = (Cg8775 | Dba775);
assign Mkg775 = (Vlg775 | H20775);
assign H20775 = (!Ht8775);
assign Ht8775 = (~(hready_i & Cmg775));
assign Cmg775 = (~(Jmg775 & Qmg775));
assign Qmg775 = (Xmg775 & Eng775);
assign Eng775 = (Lng775 & Sng775);
assign Lng775 = (~(Zng775 & Uo9775));
assign Zng775 = (Ik0775 & Bni675);
assign Xmg775 = (Gog775 & Nog775);
assign Nog775 = (~(Lzb775 & Q91775));
assign Gog775 = (~(Uog775 & E5z675));
assign Uog775 = (~(Bpg775 & Ipg775));
assign Ipg775 = (Ppg775 & Rny675);
assign Ppg775 = (~(Wpg775 & Ib9775));
assign Wpg775 = (~(Pb9775 | Dqg775));
assign Bpg775 = (Kqg775 & Rqg775);
assign Rqg775 = (~(Yqg775 & Joi675));
assign Kqg775 = (~(C1g775 & Frg775));
assign Jmg775 = (Mrg775 & Trg775);
assign Trg775 = (Asg775 & Hsg775);
assign Hsg775 = (~(Tte775 & Osg775));
assign Asg775 = (~(Mdg775 & Vsg775));
assign Mrg775 = (Ctg775 & O5b775);
assign Ctg775 = (!Jtg775);
assign Jtg775 = (Ezo675 ? Qtg775 : Jh0775);
assign Qtg775 = (Os9775 & U50775);
assign T2s675 = (Hph675 ? Eug775 : Xtg775);
assign Eug775 = (~(Lug775 & Sug775));
assign Sug775 = (Zug775 & Gvg775);
assign Zug775 = (~(Zry675 | Nvg775));
assign Lug775 = (~(Uvg775 | Bwg775));
assign Xtg775 = (~(Iwg775 & Pwg775));
assign Pwg775 = (Wwg775 & Scz675);
assign Wwg775 = (~(rxev_i | txev_o));
assign txev_o = (Dxg775 & Kxg775);
assign Dxg775 = (~(Rxg775 | Pw9775));
assign Iwg775 = (Yxg775 & Cbz675);
assign Cbz675 = (!Bt5775);
assign Bt5775 = (Fyg775 & Gtb775);
assign Yxg775 = (~(Nbp675 & Myg775));
assign Myg775 = (~(Tyg775 & Azg775));
assign Azg775 = (Hzg775 & Ozg775);
assign Ozg775 = (Vzg775 & C0h775);
assign C0h775 = (J0h775 & Q0h775);
assign Q0h775 = (X0h775 & E1h775);
assign E1h775 = (Ub8775 | E7r675);
assign Ub8775 = (L1h775 & S1h775);
assign S1h775 = (~(Z1h775 & G2h775));
assign G2h775 = (F4r675 & V72l85[0]);
assign Z1h775 = (Dg5775 & Yn5775);
assign Yn5775 = (!Wf5775);
assign Wf5775 = (~(N2h775 & U2h775));
assign U2h775 = (B3h775 & I3h775);
assign I3h775 = (P3h775 & W3h775);
assign W3h775 = (~(D4h775 | V72l85[7]));
assign D4h775 = (V72l85[8] | V72l85[9]);
assign P3h775 = (~(K4h775 | V72l85[4]));
assign K4h775 = (V72l85[5] | V72l85[6]);
assign B3h775 = (R4h775 & Y4h775);
assign Y4h775 = (~(F5h775 | V72l85[23]));
assign F5h775 = (V72l85[2] | V72l85[3]);
assign R4h775 = (~(M5h775 | V72l85[20]));
assign M5h775 = (V72l85[21] | V72l85[22]);
assign N2h775 = (T5h775 & A6h775);
assign A6h775 = (H6h775 & O6h775);
assign O6h775 = (~(V6h775 | V72l85[18]));
assign V6h775 = (V72l85[19] | V72l85[1]);
assign H6h775 = (~(C7h775 | V72l85[15]));
assign C7h775 = (V72l85[16] | V72l85[17]);
assign T5h775 = (J7h775 & Q7h775);
assign Q7h775 = (~(X7h775 | V72l85[12]));
assign X7h775 = (V72l85[13] | V72l85[14]);
assign J7h775 = (~(V72l85[10] | V72l85[11]));
assign Dg5775 = (S5r675 & E8h775);
assign E8h775 = (st_clk_en_i | L8h775);
assign L1h775 = (~(Pe6775 & hwdata_o[26]));
assign X0h775 = (S8h775 & Z8h775);
assign Z8h775 = (~(G9h775 & P58775));
assign G9h775 = (~(D68775 | Ogp675));
assign D68775 = (N9h775 & U9h775);
assign U9h775 = (~(Bah775 & Z8a775));
assign Bah775 = (Iah775 & T5a775);
assign S8h775 = (~(Pah775 & Pe6775));
assign Pah775 = (~(Uu3775 | Ifp675));
assign J0h775 = (Wah775 & Dbh775);
assign Dbh775 = (H27775 | Cep675);
assign H27775 = (Kbh775 & Rbh775);
assign Rbh775 = (N9h775 | P58775);
assign N9h775 = (~(Ybh775 & Fch775));
assign Fch775 = (~(Lrh675 | N0p675));
assign Ybh775 = (~(Mch775 | L2g775));
assign Kbh775 = (Tch775 & Adh775);
assign Adh775 = (~(Hdh775 & Odh775));
assign Odh775 = (Vdh775 & Me8775);
assign Vdh775 = (~(Of8775 & Ceh775));
assign Of8775 = (!At1775);
assign At1775 = (~(Jeh775 & Qeh775));
assign Qeh775 = (Xeh775 & Efh775);
assign Efh775 = (~(Lfh775 & Sfh775));
assign Sfh775 = (~(Wxf775 | U50775));
assign Lfh775 = (~(E5z675 | Zfh775));
assign Xeh775 = (Lvf775 & Ggh775);
assign Jeh775 = (Ngh775 & Ugh775);
assign Ngh775 = (~(Tte775 & Xza775));
assign Tte775 = (Bhh775 & Dny675);
assign Bhh775 = (~(L2g775 | Y1z675));
assign Hdh775 = (~(M71775 | Cg8775));
assign Tch775 = (~(Ihh775 & T17775));
assign Ihh775 = (~(Phh775 & Whh775));
assign Whh775 = (Dih775 & Kih775);
assign Kih775 = (~(Rih775 & Yih775));
assign Yih775 = (~(Xuf775 | Q6b775));
assign Rih775 = (Fjh775 & Nzy675);
assign Dih775 = (~(Mjh775 & Tjh775));
assign Phh775 = (Akh775 & Hkh775);
assign Hkh775 = (~(Okh775 & V8p675));
assign Okh775 = (~(Cg8775 | Me8775));
assign Wah775 = (~(Amp675 & Vkh775));
assign Vkh775 = (!Gi2l85[0]);
assign Amp675 = (R8z675 & Clh775);
assign Clh775 = (~(Jlh775 & Qlh775));
assign Qlh775 = (~(irq_i[0] & K8z675));
assign K8z675 = (!Qj2l85[0]);
assign Jlh775 = (Xlh775 & Emh775);
assign Emh775 = (~(Gi2l85[0] & Lmh775));
assign Lmh775 = (~(hwdata_o[0] & Smh775));
assign Xlh775 = (Vaz675 | Zmh775);
assign Vaz675 = (!hwdata_o[0]);
assign R8z675 = (Jbz675 | Scz675);
assign Jbz675 = (!T9z675);
assign Vzg775 = (Gnh775 & Nnh775);
assign Nnh775 = (Unh775 & Boh775);
assign Boh775 = (~(A5q675 & Ioh775));
assign Ioh775 = (!Gi2l85[12]);
assign A5q675 = (Bd7775 & Poh775);
assign Poh775 = (~(Woh775 & Dph775));
assign Dph775 = (~(irq_i[12] & Uc7775));
assign Uc7775 = (!Qj2l85[12]);
assign Woh775 = (Kph775 & Rph775);
assign Rph775 = (~(Gi2l85[12] & Yph775));
assign Yph775 = (~(Smh775 & hwdata_o[12]));
assign Kph775 = (Zmh775 | Fb4775);
assign Fb4775 = (!hwdata_o[12]);
assign Bd7775 = (Re7775 | Scz675);
assign Re7775 = (!Wd7775);
assign Unh775 = (Fqh775 & Mqh775);
assign Mqh775 = (~(U1q675 & Tqh775));
assign Tqh775 = (!Gi2l85[10]);
assign U1q675 = (Zi7775 & Arh775);
assign Arh775 = (~(Hrh775 & Orh775));
assign Orh775 = (~(irq_i[10] & Si7775));
assign Si7775 = (!Qj2l85[10]);
assign Hrh775 = (Vrh775 & Csh775);
assign Csh775 = (~(Gi2l85[10] & Jsh775));
assign Jsh775 = (~(Smh775 & hwdata_o[10]));
assign Vrh775 = (Zmh775 | Jd4775);
assign Jd4775 = (!hwdata_o[10]);
assign Zi7775 = (Pk7775 | Scz675);
assign Pk7775 = (!Uj7775);
assign Fqh775 = (~(K3q675 & Qsh775));
assign Qsh775 = (!Gi2l85[11]);
assign K3q675 = (Ag7775 & Xsh775);
assign Xsh775 = (~(Eth775 & Lth775));
assign Lth775 = (~(irq_i[11] & Tf7775));
assign Tf7775 = (!Qj2l85[11]);
assign Eth775 = (Sth775 & Zth775);
assign Zth775 = (~(Gi2l85[11] & Guh775));
assign Guh775 = (~(Smh775 & hwdata_o[11]));
assign Sth775 = (Zmh775 | Hc4775);
assign Ag7775 = (Qh7775 | Scz675);
assign Gnh775 = (Nuh775 & Uuh775);
assign Uuh775 = (~(Q6q675 & Bvh775));
assign Bvh775 = (!Gi2l85[13]);
assign Q6q675 = (Ca7775 & Ivh775);
assign Ivh775 = (~(Pvh775 & Wvh775));
assign Wvh775 = (~(irq_i[13] & V97775));
assign V97775 = (!Qj2l85[13]);
assign Pvh775 = (Dwh775 & Kwh775);
assign Kwh775 = (~(Gi2l85[13] & Rwh775));
assign Rwh775 = (~(Smh775 & hwdata_o[13]));
assign Dwh775 = (Zmh775 | Da4775);
assign Da4775 = (!hwdata_o[13]);
assign Ca7775 = (Sb7775 | Scz675);
assign Nuh775 = (~(G8q675 & Ywh775));
assign Ywh775 = (!Gi2l85[14]);
assign G8q675 = (K77775 & Fxh775);
assign Fxh775 = (~(Mxh775 & Txh775));
assign Txh775 = (~(irq_i[14] & D77775));
assign D77775 = (!Qj2l85[14]);
assign Mxh775 = (Ayh775 & Hyh775);
assign Hyh775 = (~(Gi2l85[14] & Oyh775));
assign Oyh775 = (~(Smh775 & hwdata_o[14]));
assign Ayh775 = (Zmh775 | B94775);
assign K77775 = (~(F87775 & Yf6775));
assign Hzg775 = (Vyh775 & Czh775);
assign Czh775 = (Jzh775 & Qzh775);
assign Qzh775 = (Xzh775 & E0i775);
assign E0i775 = (~(Cdq675 & L0i775));
assign L0i775 = (!Gi2l85[17]);
assign Cdq675 = (Lh8775 & S0i775);
assign S0i775 = (~(Z0i775 & G1i775));
assign G1i775 = (~(irq_i[17] & Eh8775));
assign Eh8775 = (!Qj2l85[17]);
assign Z0i775 = (Ni8775 & N1i775);
assign N1i775 = (~(Gi2l85[17] & U1i775));
assign U1i775 = (~(hwdata_o[17] & Smh775));
assign hwdata_o[17] = (!C64775);
assign Ni8775 = (C64775 | Zmh775);
assign Lh8775 = (Ui8775 | Scz675);
assign Xzh775 = (B2i775 & I2i775);
assign I2i775 = (~(W9q675 & P2i775));
assign P2i775 = (!Gi2l85[15]);
assign W9q675 = (L47775 & W2i775);
assign W2i775 = (~(D3i775 & K3i775));
assign K3i775 = (~(irq_i[15] & E47775));
assign E47775 = (!Qj2l85[15]);
assign D3i775 = (R3i775 & Y3i775);
assign Y3i775 = (~(Gi2l85[15] & F4i775));
assign F4i775 = (~(Smh775 & hwdata_o[15]));
assign R3i775 = (Zmh775 | Z74775);
assign L47775 = (B67775 | Scz675);
assign B2i775 = (~(Mbq675 & M4i775));
assign M4i775 = (!Gi2l85[16]);
assign Mbq675 = (Dk8775 & T4i775);
assign T4i775 = (~(A5i775 & H5i775));
assign H5i775 = (~(irq_i[16] & Wj8775));
assign Wj8775 = (!Qj2l85[16]);
assign A5i775 = (O5i775 & V5i775);
assign V5i775 = (~(Gi2l85[16] & C6i775));
assign C6i775 = (~(Smh775 & hwdata_o[16]));
assign O5i775 = (~(M9z675 & hwdata_o[16]));
assign Dk8775 = (J6i775 | Scz675);
assign J6i775 = (!Yk8775);
assign Jzh775 = (Q6i775 & X6i775);
assign X6i775 = (~(Seq675 & E7i775));
assign E7i775 = (!Gi2l85[18]);
assign Seq675 = (Nz5775 & L7i775);
assign L7i775 = (~(S7i775 & Z7i775));
assign Z7i775 = (~(irq_i[18] & Gz5775));
assign Gz5775 = (!Qj2l85[18]);
assign S7i775 = (G8i775 & N8i775);
assign N8i775 = (~(Gi2l85[18] & U8i775));
assign U8i775 = (~(Smh775 & hwdata_o[18]));
assign G8i775 = (Zmh775 | A54775);
assign Nz5775 = (D16775 | Scz675);
assign D16775 = (!I06775);
assign Q6i775 = (~(Igq675 & B9i775));
assign B9i775 = (!Gi2l85[19]);
assign Igq675 = (Vw5775 & I9i775);
assign I9i775 = (~(P9i775 & W9i775));
assign W9i775 = (~(irq_i[19] & Ow5775));
assign Ow5775 = (!Qj2l85[19]);
assign P9i775 = (Xx5775 & Dai775);
assign Dai775 = (~(Gi2l85[19] & Kai775));
assign Kai775 = (~(hwdata_o[19] & Smh775));
assign Xx5775 = (~(hwdata_o[19] & M9z675));
assign Vw5775 = (Ey5775 | Scz675);
assign Vyh775 = (Rai775 & Yai775);
assign Yai775 = (Fbi775 & Mbi775);
assign Mbi775 = (~(Pnp675 & Tbi775));
assign Tbi775 = (!Gi2l85[1]);
assign Pnp675 = (Ea8775 & Aci775);
assign Aci775 = (~(Hci775 & Oci775));
assign Oci775 = (~(irq_i[1] & X98775));
assign X98775 = (!Qj2l85[1]);
assign Hci775 = (Vci775 & Cdi775);
assign Cdi775 = (~(Gi2l85[1] & Jdi775));
assign Jdi775 = (~(hwdata_o[1] & Smh775));
assign Vci775 = (~(hwdata_o[1] & M9z675));
assign Ea8775 = (Qdi775 | Scz675);
assign Fbi775 = (~(Yhq675 & Xdi775));
assign Xdi775 = (!Gi2l85[20]);
assign Yhq675 = (Lc6775 & Eei775);
assign Eei775 = (~(Lei775 & Sei775));
assign Sei775 = (~(irq_i[20] & Ec6775));
assign Ec6775 = (!Qj2l85[20]);
assign Lei775 = (Nd6775 & Zei775);
assign Zei775 = (~(Gi2l85[20] & Gfi775));
assign Gfi775 = (~(hwdata_o[20] & Smh775));
assign Nd6775 = (~(hwdata_o[20] & M9z675));
assign Lc6775 = (Ud6775 | Scz675);
assign Rai775 = (Nfi775 & Ufi775);
assign Ufi775 = (~(Ojq675 & Bgi775));
assign Bgi775 = (!Gi2l85[21]);
assign Ojq675 = (T96775 & Igi775);
assign Igi775 = (~(Pgi775 & Wgi775));
assign Wgi775 = (~(irq_i[21] & M96775));
assign M96775 = (!Qj2l85[21]);
assign Pgi775 = (Va6775 & Dhi775);
assign Dhi775 = (~(Gi2l85[21] & Khi775));
assign Khi775 = (~(hwdata_o[21] & Smh775));
assign Va6775 = (~(hwdata_o[21] & M9z675));
assign T96775 = (Cb6775 | Scz675);
assign Nfi775 = (~(Elq675 & Rhi775));
assign Rhi775 = (!Gi2l85[22]);
assign Elq675 = (U66775 & Yhi775);
assign Yhi775 = (~(Fii775 & Mii775));
assign Mii775 = (~(irq_i[22] & N66775));
assign N66775 = (!Qj2l85[22]);
assign Fii775 = (Tii775 & Aji775);
assign Aji775 = (~(Gi2l85[22] & Hji775));
assign Hji775 = (~(Smh775 & hwdata_o[22]));
assign Tii775 = (Zmh775 | G14775);
assign U66775 = (K86775 | Scz675);
assign K86775 = (!P76775);
assign Tyg775 = (Oji775 & Vji775);
assign Vji775 = (Cki775 & Jki775);
assign Jki775 = (Qki775 & Xki775);
assign Xki775 = (Eli775 & Lli775);
assign Lli775 = (~(Aqq675 & Sli775));
assign Aqq675 = (Yz7775 & Zli775);
assign Zli775 = (~(Gmi775 & Nmi775));
assign Nmi775 = (~(irq_i[25] & Rz7775));
assign Rz7775 = (!Qj2l85[25]);
assign Gmi775 = (Umi775 & Bni775);
assign Bni775 = (~(Gi2l85[25] & Ini775));
assign Ini775 = (~(Smh775 & hwdata_o[25]));
assign Umi775 = (Zmh775 | Ay3775);
assign Ay3775 = (!hwdata_o[25]);
assign Yz7775 = (O18775 | Scz675);
assign Eli775 = (Pni775 & Wni775);
assign Wni775 = (~(Umq675 & Doi775));
assign Doi775 = (!Gi2l85[23]);
assign Umq675 = (C46775 & Koi775);
assign Koi775 = (~(Roi775 & Yoi775));
assign Yoi775 = (~(irq_i[23] & V36775));
assign V36775 = (!Qj2l85[23]);
assign Roi775 = (E56775 & Fpi775);
assign Fpi775 = (~(Gi2l85[23] & Mpi775));
assign Mpi775 = (~(hwdata_o[23] & Smh775));
assign E56775 = (E04775 | Zmh775);
assign C46775 = (L56775 | Scz675);
assign Pni775 = (~(Koq675 & Tpi775));
assign Tpi775 = (!Gi2l85[24]);
assign Koq675 = (X28775 & Aqi775);
assign Aqi775 = (~(Hqi775 & Oqi775));
assign Oqi775 = (~(irq_i[24] & Q28775));
assign Q28775 = (!Qj2l85[24]);
assign Hqi775 = (Z38775 & Vqi775);
assign Vqi775 = (~(Gi2l85[24] & Cri775));
assign Cri775 = (~(Smh775 & hwdata_o[24]));
assign Z38775 = (Zmh775 | Cz3775);
assign X28775 = (G48775 | Scz675);
assign G48775 = (!Jri775);
assign Qki775 = (Qri775 & Xri775);
assign Xri775 = (~(Qrq675 & Esi775));
assign Esi775 = (!Gi2l85[26]);
assign Qrq675 = (Gx7775 & Lsi775);
assign Lsi775 = (~(Ssi775 & Zsi775));
assign Zsi775 = (~(irq_i[26] & Zw7775));
assign Zw7775 = (!Qj2l85[26]);
assign Ssi775 = (Iy7775 & Gti775);
assign Gti775 = (~(Gi2l85[26] & Nti775));
assign Nti775 = (~(Smh775 & hwdata_o[26]));
assign Iy7775 = (Zmh775 | Yw3775);
assign Gx7775 = (Py7775 | Scz675);
assign Py7775 = (!Uti775);
assign Qri775 = (~(Gtq675 & Bui775));
assign Gtq675 = (Hu7775 & Iui775);
assign Iui775 = (~(Pui775 & Wui775));
assign Wui775 = (~(irq_i[27] & Au7775));
assign Au7775 = (!Qj2l85[27]);
assign Pui775 = (Dvi775 & Kvi775);
assign Kvi775 = (~(Gi2l85[27] & Rvi775));
assign Rvi775 = (~(Smh775 & hwdata_o[27]));
assign Dvi775 = (Zmh775 | Wv3775);
assign Wv3775 = (!hwdata_o[27]);
assign Hu7775 = (Xv7775 | Scz675);
assign Cki775 = (Yvi775 & Fwi775);
assign Fwi775 = (Mwi775 & Twi775);
assign Twi775 = (~(Wuq675 & Axi775));
assign Axi775 = (!Gi2l85[28]);
assign Wuq675 = (Pr7775 & Hxi775);
assign Hxi775 = (~(Oxi775 & Vxi775));
assign Vxi775 = (~(irq_i[28] & Ir7775));
assign Ir7775 = (!Qj2l85[28]);
assign Oxi775 = (Rs7775 & Cyi775);
assign Cyi775 = (~(Gi2l85[28] & Jyi775));
assign Jyi775 = (~(Smh775 & hwdata_o[28]));
assign Rs7775 = (Zmh775 | Uu3775);
assign Uu3775 = (!hwdata_o[28]);
assign Pr7775 = (Ys7775 | Scz675);
assign Ys7775 = (!Qyi775);
assign Mwi775 = (~(Mwq675 & Xyi775));
assign Mwq675 = (Gs5775 & Ezi775);
assign Ezi775 = (~(Lzi775 & Szi775));
assign Szi775 = (~(irq_i[29] & Zr5775));
assign Zr5775 = (!Qj2l85[29]);
assign Lzi775 = (Pt5775 & Zzi775);
assign Zzi775 = (~(Gi2l85[29] & G0j775));
assign G0j775 = (~(Smh775 & hwdata_o[29]));
assign Pt5775 = (Zmh775 | St3775);
assign St3775 = (!hwdata_o[29]);
assign Gs5775 = (Wt5775 | Scz675);
assign Yvi775 = (N0j775 & U0j775);
assign U0j775 = (~(Epp675 & B1j775));
assign B1j775 = (!Gi2l85[2]);
assign Epp675 = (M78775 & I1j775);
assign I1j775 = (~(P1j775 & W1j775));
assign W1j775 = (~(irq_i[2] & F78775));
assign F78775 = (!Qj2l85[2]);
assign P1j775 = (O88775 & D2j775);
assign D2j775 = (~(Gi2l85[2] & K2j775));
assign K2j775 = (~(Xk4775 & Smh775));
assign O88775 = (~(Xk4775 & M9z675));
assign M78775 = (V88775 | Scz675);
assign N0j775 = (~(Cyq675 & R2j775));
assign R2j775 = (!Gi2l85[30]);
assign Cyq675 = (Vm8775 & Y2j775);
assign Y2j775 = (~(F3j775 & M3j775));
assign M3j775 = (~(irq_i[30] & Om8775));
assign Om8775 = (!Qj2l85[30]);
assign F3j775 = (T3j775 & A4j775);
assign A4j775 = (~(Gi2l85[30] & H4j775));
assign H4j775 = (~(Smh775 & hwdata_o[30]));
assign T3j775 = (Zmh775 | Qs3775);
assign Qs3775 = (!hwdata_o[30]);
assign Vm8775 = (Lo8775 | Scz675);
assign Lo8775 = (!Qn8775);
assign Oji775 = (O4j775 & V4j775);
assign V4j775 = (C5j775 & J5j775);
assign J5j775 = (Q5j775 & X5j775);
assign X5j775 = (~(Isp675 & E6j775));
assign E6j775 = (!Gi2l85[4]);
assign Isp675 = (Gr6775 & L6j775);
assign L6j775 = (~(S6j775 & Z6j775));
assign Z6j775 = (~(irq_i[4] & Zq6775));
assign Zq6775 = (!Qj2l85[4]);
assign S6j775 = (G7j775 & N7j775);
assign N7j775 = (~(Gi2l85[4] & U7j775));
assign U7j775 = (~(hwdata_o[4] & Smh775));
assign G7j775 = (Aj4775 | Zmh775);
assign Aj4775 = (!hwdata_o[4]);
assign Gr6775 = (Ws6775 | Scz675);
assign Ws6775 = (!Bs6775);
assign Q5j775 = (B8j775 & I8j775);
assign I8j775 = (~(Szq675 & P8j775));
assign P8j775 = (!Gi2l85[31]);
assign Szq675 = (Hp5775 & W8j775);
assign W8j775 = (~(D9j775 & K9j775));
assign K9j775 = (~(irq_i[31] & Ap5775));
assign Ap5775 = (!Qj2l85[31]);
assign D9j775 = (R9j775 & Y9j775);
assign Y9j775 = (~(Gi2l85[31] & Faj775));
assign Faj775 = (~(Smh775 & hwdata_o[31]));
assign R9j775 = (Zmh775 | Nyz675);
assign Hp5775 = (Xq5775 | Scz675);
assign B8j775 = (~(Tqp675 & Maj775));
assign Maj775 = (!Gi2l85[3]);
assign Tqp675 = (Fu6775 & Taj775);
assign Taj775 = (~(Abj775 & Hbj775));
assign Hbj775 = (~(irq_i[3] & Yt6775));
assign Yt6775 = (!Qj2l85[3]);
assign Abj775 = (Obj775 & Vbj775);
assign Vbj775 = (~(Gi2l85[3] & Ccj775));
assign Ccj775 = (~(hwdata_o[3] & Smh775));
assign Obj775 = (~(hwdata_o[3] & M9z675));
assign Fu6775 = (Jcj775 | Scz675);
assign C5j775 = (Qcj775 & Xcj775);
assign Xcj775 = (~(Xtp675 & Edj775));
assign Edj775 = (!Gi2l85[5]);
assign Xtp675 = (Ho6775 & Ldj775);
assign Ldj775 = (~(Sdj775 & Zdj775));
assign Zdj775 = (~(irq_i[5] & Ao6775));
assign Ao6775 = (!Qj2l85[5]);
assign Sdj775 = (Gej775 & Nej775);
assign Nej775 = (~(Gi2l85[5] & Uej775));
assign Uej775 = (~(hwdata_o[5] & Smh775));
assign Gej775 = (Yh4775 | Zmh775);
assign Yh4775 = (!hwdata_o[5]);
assign Ho6775 = (Xp6775 | Scz675);
assign Qcj775 = (~(Mvp675 & Bfj775));
assign Bfj775 = (!Gi2l85[6]);
assign Mvp675 = (Pl6775 & Ifj775);
assign Ifj775 = (~(Pfj775 & Wfj775));
assign Wfj775 = (~(irq_i[6] & Il6775));
assign Il6775 = (!Qj2l85[6]);
assign Pfj775 = (Dgj775 & Kgj775);
assign Kgj775 = (~(Gi2l85[6] & Rgj775));
assign Rgj775 = (~(hwdata_o[6] & Smh775));
assign Dgj775 = (~(hwdata_o[6] & M9z675));
assign Pl6775 = (Ygj775 | Scz675);
assign Ygj775 = (!Km6775);
assign O4j775 = (Fhj775 & Mhj775);
assign Mhj775 = (Thj775 & Aij775);
assign Aij775 = (~(Bxp675 & Hij775));
assign Hij775 = (!Gi2l85[7]);
assign Bxp675 = (Xi6775 & Oij775);
assign Oij775 = (~(Vij775 & Cjj775));
assign Cjj775 = (~(irq_i[7] & Qi6775));
assign Qi6775 = (!Qj2l85[7]);
assign Vij775 = (Jjj775 & Qjj775);
assign Qjj775 = (~(Gi2l85[7] & Xjj775));
assign Xjj775 = (~(hwdata_o[7] & Smh775));
assign Jjj775 = (~(hwdata_o[7] & M9z675));
assign Xi6775 = (Ekj775 | Scz675);
assign Thj775 = (~(Qyp675 & Lkj775));
assign Lkj775 = (!Gi2l85[8]);
assign Qyp675 = (Qo7775 & Skj775);
assign Skj775 = (~(Zkj775 & Glj775));
assign Glj775 = (~(irq_i[8] & Jo7775));
assign Jo7775 = (!Qj2l85[8]);
assign Zkj775 = (Nlj775 & Ulj775);
assign Ulj775 = (~(Gi2l85[8] & Bmj775));
assign Bmj775 = (~(Smh775 & hwdata_o[8]));
assign Nlj775 = (Zmh775 | Gf4775);
assign Qo7775 = (Gq7775 | Scz675);
assign Fhj775 = (Imj775 & Pmj775);
assign Pmj775 = (~(F0q675 & Wmj775));
assign Wmj775 = (!Gi2l85[9]);
assign F0q675 = (Yl7775 & Dnj775);
assign Dnj775 = (~(Knj775 & Rnj775));
assign Rnj775 = (~(irq_i[9] & Rl7775));
assign Rl7775 = (!Qj2l85[9]);
assign Knj775 = (Ynj775 & Foj775);
assign Foj775 = (~(Gi2l85[9] & Moj775));
assign Moj775 = (~(Smh775 & hwdata_o[9]));
assign Smh775 = (Gm4775 & Toj775);
assign Gm4775 = (~(Or3775 | Apj775));
assign Or3775 = (!Lnh675);
assign Ynj775 = (~(M9z675 & hwdata_o[9]));
assign M9z675 = (!Zmh775);
assign Zmh775 = (~(Hpj775 & Opj775));
assign Hpj775 = (Toj775 & Lnh675);
assign Yl7775 = (~(Tm7775 & Yf6775));
assign Yf6775 = (!Scz675);
assign Imj775 = (~(Gjp675 & Vpj775));
assign Gjp675 = (Pz6775 & Cqj775);
assign Cqj775 = (~(Jqj775 & Qqj775));
assign Qqj775 = (~(nmi_i & Iz6775));
assign Iz6775 = (!Skp675);
assign Jqj775 = (Bz6775 & Vpj775);
assign Bz6775 = (~(Pe6775 & hwdata_o[31]));
assign Pe6775 = (Lnh675 & Xqj775);
assign Pz6775 = (Scz675 | D07775);
assign D07775 = (!Erj775);
assign Scz675 = (~(Lrj775 & Srj775));
assign Lrj775 = (Zrj775 & Sfa775);
assign Sfa775 = (~(U50775 | Lrh675));
assign Y1s675 = (!Gsj775);
assign Gsj775 = (hready_i ? Usj775 : Nsj775);
assign Usj775 = (Btj775 & Itj775);
assign Itj775 = (Ptj775 & Wtj775);
assign Wtj775 = (Duj775 & Kuj775);
assign Kuj775 = (~(Ruj775 & Yuj775));
assign Ruj775 = (Fvj775 & Hk3775);
assign Fvj775 = (Mvj775 | Gw8775);
assign Duj775 = (Tvj775 & Awj775);
assign Awj775 = (~(Hwj775 & Owj775));
assign Hwj775 = (Vwj775 & Cxj775);
assign Cxj775 = (~(Iq1775 ^ Jxj775));
assign Tvj775 = (~(Qxj775 & Xxj775));
assign Qxj775 = (Bni675 & Eyj775);
assign Eyj775 = (Lyj775 | Tc3775);
assign Ptj775 = (Syj775 & Zyj775);
assign Zyj775 = (~(Gzj775 & Osg775));
assign Gzj775 = (~(Ibg775 | Mwo675));
assign Syj775 = (~(Gtb775 & Nzj775));
assign Nzj775 = (~(Uzj775 & B0k775));
assign B0k775 = (~(I0k775 & Dba775));
assign I0k775 = (Dny675 & X7a775);
assign Uzj775 = (Ep0775 | Rto675);
assign Btj775 = (P0k775 & W0k775);
assign W0k775 = (D1k775 & K1k775);
assign K1k775 = (~(Wk0775 & C1g775));
assign D1k775 = (R1k775 & Y1k775);
assign Y1k775 = (~(Ub1775 & F2k775));
assign F2k775 = (~(M2k775 & T2k775));
assign T2k775 = (~(A3k775 & Sh1775));
assign R1k775 = (~(F6g775 & H3k775));
assign H3k775 = (~(O3k775 & V3k775));
assign V3k775 = (~(Osg775 & C4k775));
assign C4k775 = (~(Rba775 & J4k775));
assign J4k775 = (O6a775 | Lrh675);
assign P0k775 = (~(Q4k775 | X4k775));
assign R1s675 = (E5k775 & L5k775);
assign L5k775 = (~(S5k775 & Z5k775));
assign Z5k775 = (G6k775 & N6k775);
assign N6k775 = (U6k775 & B7k775);
assign B7k775 = (Wub775 & Ggh775);
assign U6k775 = (I7k775 & P7k775);
assign P7k775 = (~(W7k775 & D8k775));
assign D8k775 = (~(U50775 | O6a775));
assign W7k775 = (~(Fkg775 | D1z675));
assign I7k775 = (~(K8k775 & Os9775));
assign K8k775 = (~(X7a775 | Ezo675));
assign G6k775 = (R8k775 & Y8k775);
assign Y8k775 = (~(F9k775 & M71775));
assign F9k775 = (~(M9k775 & T9k775));
assign T9k775 = (Aak775 & Hak775);
assign Hak775 = (~(Oak775 & Kq9775));
assign Oak775 = (~(Pb9775 | Gwh675));
assign Aak775 = (Vak775 & C7a775);
assign C7a775 = (~(Cbk775 & D3b775));
assign Cbk775 = (~(Jbk775 | X5p675));
assign M9k775 = (Qbk775 & Xbk775);
assign Xbk775 = (~(Zx6775 & Frg775));
assign Qbk775 = (~(Eck775 & Zfa775));
assign R8k775 = (Lck775 & Sck775);
assign Sck775 = (~(Zck775 & Gdk775));
assign Gdk775 = (~(Ndk775 & Udk775));
assign Udk775 = (~(My9775 & Bek775));
assign Lck775 = (~(Iek775 & Pek775));
assign Pek775 = (~(Wek775 & Dfk775));
assign Dfk775 = (~(Kfk775 & Rfk775));
assign Rfk775 = (Yfk775 & Fgk775);
assign Kfk775 = (Mgk775 & Tgk775);
assign Mgk775 = (~(Nh9775 | Ahk775));
assign Wek775 = (~(Hhk775 | Bk0775));
assign S5k775 = (Ohk775 & Vhk775);
assign Vhk775 = (Cik775 & Jik775);
assign Cik775 = (Qik775 & Xik775);
assign Xik775 = (~(Gwf775 & Ejk775));
assign Ejk775 = (~(Ljk775 & Sjk775));
assign Sjk775 = (~(Ib9775 & Zjk775));
assign Zjk775 = (~(Gkk775 & Nkk775));
assign Nkk775 = (~(Lki675 | Bni675));
assign Gkk775 = (Ukk775 & Blk775);
assign Blk775 = (~(Ilk775 ^ Eji675));
assign Ukk775 = (M53775 ? Qgi675 : Lyj775);
assign Ljk775 = (Plk775 & Wlk775);
assign Wlk775 = (~(O79775 & Dmk775));
assign Dmk775 = (~(Ye0775 & Kmk775));
assign Kmk775 = (Tc3775 | Ef3775);
assign Plk775 = (~(Zqi675 & Rmk775));
assign Rmk775 = (~(Ymk775 & Fnk775));
assign Fnk775 = (~(Mnk775 & Hk3775));
assign Mnk775 = (~(Tnk775 & Aok775));
assign Aok775 = (Tli675 ? Ook775 : Hok775);
assign Ook775 = (~(Vok775 & Cpk775));
assign Cpk775 = (~(Ia3775 | M53775));
assign Vok775 = (Jpk775 & Qpk775);
assign Hok775 = (!Xpk775);
assign Tnk775 = (Joi675 & Eqk775);
assign Ymk775 = (~(Lqk775 & Sqk775));
assign Sqk775 = (~(M53775 ^ Zqk775));
assign Lqk775 = (~(Dc9775 | Joi675));
assign Qik775 = (B2b775 | Za1775);
assign Ohk775 = (~(Grk775 | Nrk775));
assign Nrk775 = (Hk3775 ? Bsk775 : Urk775);
assign Urk775 = (Hs9775 & Ria775);
assign Hs9775 = (Isk775 & Uag775);
assign Isk775 = (Jf9775 & Psk775);
assign Grk775 = (Wsk775 | Dtk775);
assign E5k775 = (Gvo675 | hready_i);
assign K1s675 = (!Ktk775);
assign Ktk775 = (hready_i ? Rtk775 : Cm2775);
assign Rtk775 = (Ytk775 & Fuk775);
assign Fuk775 = (Muk775 & Tuk775);
assign Tuk775 = (Avk775 & Hvk775);
assign Hvk775 = (Ovk775 & Vvk775);
assign Vvk775 = (~(Cwk775 & Jwk775));
assign Jwk775 = (Qwk775 & Rj9775);
assign Qwk775 = (~(Dc9775 | V8p675));
assign Cwk775 = (Xwk775 & Ik0775);
assign Xwk775 = (Zqk775 ^ M53775);
assign Zqk775 = (Exk775 & Lxk775);
assign Lxk775 = (Sxk775 ^ Zxk775);
assign Zxk775 = (Gyk775 & Nyk775);
assign Nyk775 = (~(Xv0775 | Owj775));
assign Xv0775 = (vis_apsr_o[0] & Gx0775);
assign Gyk775 = (Uyk775 & Bzk775);
assign Bzk775 = (Tli675 | Izk775);
assign Uyk775 = (Pzk775 | Wzk775);
assign Wzk775 = (Kq1l85 ? Sy1l85[31] : Rjl675);
assign Pzk775 = (D0l775 | Gx0775);
assign Gx0775 = (K0l775 & R0l775);
assign K0l775 = (Y0l775 & F1l775);
assign F1l775 = (~(M1l775 & T1l775));
assign T1l775 = (~(Pw9775 | Xza775));
assign M1l775 = (~(A2l775 | Veg775));
assign Y0l775 = (~(H2l775 & Rcg775));
assign H2l775 = (~(O2l775 | Cm2775));
assign D0l775 = (~(Rjl675 | Sy1l85[31]));
assign Rjl675 = (~(V2l775 | Foy675));
assign Foy675 = (!Jqy675);
assign Jqy675 = (~(C3l775 & J3l775));
assign J3l775 = (Q3l775 & X3l775);
assign X3l775 = (E4l775 & L4l775);
assign L4l775 = (Bwg775 | Bbg775);
assign E4l775 = (Xuf775 | X5p675);
assign Q3l775 = (S4l775 & Z4l775);
assign Z4l775 = (Yyf775 | Y1z675);
assign S4l775 = (Te1775 | Q91775);
assign C3l775 = (G5l775 & N5l775);
assign N5l775 = (N0p675 ? B6l775 : U5l775);
assign B6l775 = (I6l775 | Q6b775);
assign U5l775 = (P6l775 & W6l775);
assign W6l775 = (U50775 | X5p675);
assign P6l775 = (~(D7l775 | Vxo675));
assign G5l775 = (K7l775 & Gvo675);
assign K7l775 = (Xza775 ? B0z675 : Rxg775);
assign Sxk775 = (R7l775 | Y7l775);
assign Y7l775 = (Sgg775 ? vis_apsr_o[3] : Iig775);
assign Iig775 = (!F8l775);
assign F8l775 = (C4i675 ? M8l775 : I1c775);
assign R7l775 = (~(T8l775 & A9l775));
assign T8l775 = (X73775 | Tli675);
assign Exk775 = (H9l775 & O9l775);
assign O9l775 = (V9l775 | Cal775);
assign Cal775 = (Uq0775 ? vis_apsr_o[1] : Rs0775);
assign Uq0775 = (Jal775 & R0l775);
assign R0l775 = (Qal775 & Xal775);
assign Xal775 = (~(Bvh675 & Ebl775));
assign Ebl775 = (~(Lbl775 & Sbl775));
assign Lbl775 = (~(Zbl775 & Kny675));
assign Zbl775 = (~(N0p675 | O4p675));
assign Qal775 = (Gcl775 & Ncl775);
assign Jal775 = (Ucl775 & Bdl775);
assign Bdl775 = (~(Bvh675 & Idl775));
assign Idl775 = (~(Pdl775 & Wdl775));
assign Pdl775 = (Del775 | O4p675);
assign Ucl775 = (~(N0p675 & Kel775));
assign Kel775 = (~(Rel775 & Yel775));
assign Yel775 = (Y1z675 | O4p675);
assign Rel775 = (Ffl775 & Mfl775);
assign Mfl775 = (~(M6g775 & Tfl775));
assign Tfl775 = (Zry675 | F6g775);
assign Ffl775 = (Agl775 | Veg775);
assign Rs0775 = (C4i675 ? Hgl775 : F6j675);
assign Hgl775 = (Vgl775 ? vis_apsr_o[1] : Ogl775);
assign Vgl775 = (Chl775 & Jhl775);
assign Chl775 = (Qhl775 & Xhl775);
assign Ogl775 = (~(Eil775 & Lil775));
assign Lil775 = (~(Sil775 & Zil775));
assign Zil775 = (~(Gjl775 & Njl775));
assign Njl775 = (Ujl775 & Bkl775);
assign Bkl775 = (Ikl775 | Pkl775);
assign Ikl775 = (Kll775 ? Dll775 : Wkl775);
assign Ujl775 = (Rll775 | Yll775);
assign Gjl775 = (Fml775 & Mml775);
assign Mml775 = (Tml775 | Anl775);
assign Fml775 = (Hnl775 | Onl775);
assign Sil775 = (Vnl775 ? Y1z675 : Zry675);
assign Eil775 = (Vnl775 ? Jol775 : Col775);
assign Vnl775 = (Xhl775 & Qol775);
assign Qol775 = (Qhl775 | Jhl775);
assign Jol775 = (~(Rto675 & Xol775));
assign Xol775 = (~(Epl775 & Lpl775));
assign Lpl775 = (Spl775 & Zpl775);
assign Zpl775 = (Gql775 | Tml775);
assign Spl775 = (Nql775 | Rll775);
assign Epl775 = (Uql775 & Brl775);
assign Brl775 = (Irl775 | Onl775);
assign Uql775 = (Prl775 | Pkl775);
assign Col775 = (M8l775 | Wrl775);
assign M8l775 = (Dsl775 & Ksl775);
assign Ksl775 = (Rsl775 & Ysl775);
assign Ysl775 = (~(Ftl775 & Mtl775));
assign Ftl775 = (~(Ttl775 & Aul775));
assign Aul775 = (Hnl775 | Hul775);
assign Ttl775 = (Oul775 | Yll775);
assign Rsl775 = (Vul775 | Cvl775);
assign Vul775 = (!Jvl775);
assign Dsl775 = (Qvl775 & Xvl775);
assign Xvl775 = (Ewl775 | Lwl775);
assign Qvl775 = (Swl775 | Anl775);
assign V9l775 = (~(Zwl775 & Ia3775));
assign Zwl775 = (~(X73775 ^ Tli675));
assign H9l775 = (~(Gxl775 & Nxl775));
assign Nxl775 = (~(Uxl775 & A9l775));
assign Uxl775 = (Tc3775 | Eji675);
assign Gxl775 = (Dqg775 ^ Byl775);
assign Byl775 = (Sgg775 ? vis_apsr_o[2] : S6c775);
assign Sgg775 = (Iyl775 & Evf775);
assign Evf775 = (Pyl775 | Veg775);
assign Iyl775 = (~(Bvh675 & Wyl775));
assign Wyl775 = (~(Dzl775 & Kzl775));
assign Kzl775 = (Rzl775 & Yzl775);
assign Yzl775 = (~(F0m775 & D1z675));
assign F0m775 = (~(M0m775 & Ezo675));
assign M0m775 = (~(T0m775 | Rto675));
assign Rzl775 = (A1m775 & Sbl775);
assign Sbl775 = (~(H1m775 & Rto675));
assign H1m775 = (O1m775 & V1m775);
assign O1m775 = (Bbg775 | Pw9775);
assign A1m775 = (V1m775 | Pw9775);
assign Dzl775 = (C2m775 & J2m775);
assign J2m775 = (Nvg775 | F3p675);
assign C2m775 = (~(Rcg775 & Kny675));
assign S6c775 = (!Q2m775);
assign Q2m775 = (C4i675 ? E3m775 : X2m775);
assign E3m775 = (~(L3m775 & S3m775));
assign S3m775 = (Z3m775 & G4m775);
assign G4m775 = (~(N4m775 & U4m775));
assign U4m775 = (Mtl775 | B5m775);
assign N4m775 = (I5m775 & P5m775);
assign I5m775 = (~(W5m775 & D6m775));
assign D6m775 = (K6m775 & R6m775);
assign K6m775 = (Yll775 & Irl775);
assign W5m775 = (Y6m775 & F7m775);
assign Y6m775 = (Kll775 ? T7m775 : M7m775);
assign T7m775 = (A8m775 & H8m775);
assign H8m775 = (O8m775 & V8m775);
assign A8m775 = (~(C9m775 | J9m775));
assign M7m775 = (Q9m775 & X9m775);
assign X9m775 = (Eam775 & Lam775);
assign Z3m775 = (Sam775 & Zam775);
assign Zam775 = (~(Gbm775 & Nbm775));
assign Nbm775 = (Ubm775 | B5m775);
assign Gbm775 = (Bcm775 & P5m775);
assign Bcm775 = (~(Icm775 & Pcm775));
assign Pcm775 = (Wcm775 & Ddm775);
assign Wcm775 = (Anl775 & Nql775);
assign Icm775 = (Kdm775 & Rdm775);
assign Kdm775 = (Kll775 ? Fem775 : Ydm775);
assign Fem775 = (Mem775 & Tem775);
assign Tem775 = (Afm775 & Hfm775);
assign Afm775 = (!Ofm775);
assign Mem775 = (Vfm775 & Cgm775);
assign Cgm775 = (!Jgm775);
assign Ydm775 = (Qgm775 & Xgm775);
assign Xgm775 = (O8m775 & Ehm775);
assign Qgm775 = (~(Lhm775 | J9m775));
assign Sam775 = (~(Shm775 & Zhm775));
assign Zhm775 = (Gim775 | Nim775);
assign L3m775 = (Uim775 & Bjm775);
assign Bjm775 = (~(Ijm775 & Pjm775));
assign Pjm775 = (~(Wjm775 & Dkm775));
assign Dkm775 = (~(Kkm775 | Rkm775));
assign Wjm775 = (Onl775 & Rll775);
assign Ijm775 = (Ykm775 & Flm775);
assign Ykm775 = (~(Mlm775 & Tlm775));
assign Tlm775 = (Amm775 & Hmm775);
assign Hmm775 = (Omm775 & Vmm775);
assign Omm775 = (Cnm775 & Jnm775);
assign Amm775 = (Qnm775 & Xnm775);
assign Mlm775 = (Eom775 & Lom775);
assign Lom775 = (Som775 & Zom775);
assign Zom775 = (~(Gpm775 & Npm775));
assign Som775 = (Upm775 & Bqm775);
assign Upm775 = (~(Iqm775 & Pqm775));
assign Pqm775 = (Wqm775 | Gpm775);
assign Eom775 = (Cvl775 & Drm775);
assign Drm775 = (~(Wqm775 & Krm775));
assign Uim775 = (~(Rrm775 & Yrm775));
assign Yrm775 = (~(Fsm775 & Msm775));
assign Msm775 = (Tsm775 & Atm775);
assign Tsm775 = (Hnl775 & Prl775);
assign Fsm775 = (Htm775 & Otm775);
assign Htm775 = (Kll775 ? Cum775 : Vtm775);
assign Cum775 = (Q9m775 & Jum775);
assign Jum775 = (Qum775 & Xum775);
assign Q9m775 = (~(Evm775 | Lvm775));
assign Vtm775 = (Svm775 & Zvm775);
assign Zvm775 = (Dll775 & Gwm775);
assign Svm775 = (~(Npm775 | Krm775));
assign Rrm775 = (~(Nwm775 & Uwm775));
assign Nwm775 = (Bxm775 & Swl775);
assign X2m775 = (~(Ixm775 & Pxm775));
assign Pxm775 = (Wxm775 & Dym775);
assign Dym775 = (Kym775 & Rym775);
assign Rym775 = (Yym775 & Fzm775);
assign Fzm775 = (Mzm775 & Tzm775);
assign Tzm775 = (~(Tz1l85[6] | Tz1l85[8]));
assign Mzm775 = (~(Tz1l85[25] | Tz1l85[26]));
assign Yym775 = (~(A0n775 | Tz1l85[20]));
assign A0n775 = (Tz1l85[21] | Tz1l85[22]);
assign Kym775 = (H0n775 & O0n775);
assign O0n775 = (V0n775 & Hvd775);
assign Hvd775 = (!Tz1l85[17]);
assign V0n775 = (~(Tz1l85[18] | Tz1l85[19]));
assign H0n775 = (~(C1n775 | Tz1l85[14]));
assign C1n775 = (Tz1l85[15] | Tz1l85[16]);
assign Wxm775 = (J1n775 & Q1n775);
assign Q1n775 = (X1n775 & E2n775);
assign E2n775 = (L2n775 & S2n775);
assign S2n775 = (~(Tz1l85[12] | Tz1l85[13]));
assign L2n775 = (Z2n775 & One775);
assign One775 = (!Tz1l85[11]);
assign Z2n775 = (~(Mbb775 & G3n775));
assign G3n775 = (~(N3n775 & U3n775));
assign U3n775 = (B4n775 & I4n775);
assign I4n775 = (P4n775 & W4n775);
assign W4n775 = (~(D5n775 | Sy1l85[3]));
assign D5n775 = (Sy1l85[6] | Sy1l85[8]);
assign P4n775 = (~(Sy1l85[26] | Sy1l85[30]));
assign B4n775 = (K5n775 & R5n775);
assign R5n775 = (~(Y5n775 | Sy1l85[21]));
assign Y5n775 = (Sy1l85[22] | Sy1l85[25]);
assign K5n775 = (~(Sy1l85[19] | Sy1l85[20]));
assign N3n775 = (F6n775 & M6n775);
assign M6n775 = (T6n775 & A7n775);
assign A7n775 = (~(H7n775 | Sy1l85[16]));
assign H7n775 = (Sy1l85[17] | Sy1l85[18]);
assign T6n775 = (~(Sy1l85[14] | Sy1l85[15]));
assign F6n775 = (O7n775 & V7n775);
assign V7n775 = (~(Sy1l85[12] | Sy1l85[13]));
assign O7n775 = (~(Sy1l85[0] | Sy1l85[11]));
assign X1n775 = (C8n775 & Hne775);
assign Hne775 = (~(J8n775 & Q8n775));
assign J8n775 = (Ct1l85 ? E9n775 : X8n775);
assign C8n775 = (~(U4f775 | L9n775));
assign L9n775 = (Ifc775 & S9n775);
assign S9n775 = (~(Z9n775 & Gan775));
assign Gan775 = (Nan775 & Uan775);
assign Uan775 = (Bbn775 & Ibn775);
assign Ibn775 = (Pbn775 & Wbn775);
assign Wbn775 = (~(Bty675 & As1l85));
assign Pbn775 = (Dcn775 & Kcn775);
assign Kcn775 = (~(Apy675 & Dq1l85));
assign Dcn775 = (~(Moy675 & Wp1l85));
assign Bbn775 = (Rcn775 & Ycn775);
assign Ycn775 = (~(Ity675 & Tr1l85));
assign Rcn775 = (~(Ruy675 & Bw1l85));
assign Nan775 = (Fdn775 & Mdn775);
assign Mdn775 = (Tdn775 & Aen775);
assign Aen775 = (~(Fvy675 & Gv1l85));
assign Tdn775 = (Hen775 & Oen775);
assign Oen775 = (~(Duy675 & Uv1l85));
assign Hen775 = (~(Kuy675 & Nv1l85));
assign Fdn775 = (Ven775 & Cfn775);
assign Cfn775 = (~(Mvy675 & Zu1l85));
assign Ven775 = (~(Hwy675 & Su1l85));
assign Z9n775 = (Jfn775 & Qfn775);
assign Qfn775 = (Xfn775 & Egn775);
assign Egn775 = (Lgn775 & Sgn775);
assign Sgn775 = (~(Owy675 & Xt1l85));
assign Lgn775 = (Zgn775 & Ghn775);
assign Ghn775 = (~(Tvy675 & Lu1l85));
assign Zgn775 = (~(Awy675 & Eu1l85));
assign Xfn775 = (Nhn775 & Uhn775);
assign Uhn775 = (~(Vwy675 & Qt1l85));
assign Nhn775 = (~(Cxy675 & Jt1l85));
assign Jfn775 = (Bin775 & Iin775);
assign Iin775 = (Pin775 & Win775);
assign Win775 = (Q8n775 | Qoe775);
assign Qoe775 = (!Ct1l85);
assign Ct1l85 = (~(Djn775 ^ Kjn775));
assign Djn775 = (~(Rjn775 & Yjn775));
assign Yjn775 = (~(Lki675 & Fkn775));
assign Rjn775 = (Mkn775 & Tkn775);
assign Mkn775 = (Aln775 | Xoe775);
assign Q8n775 = (!Jxy675);
assign Jxy675 = (Oln775 ? Bke775 : Hln775);
assign Bke775 = (!J0m675);
assign Hln775 = (Vln775 & Cmn775);
assign Cmn775 = (Jmn775 & Qmn775);
assign Qmn775 = (Xmn775 & Enn775);
assign Enn775 = (~(Lnn775 & vis_r14_o[11]));
assign Xmn775 = (Snn775 & Znn775);
assign Znn775 = (~(Gon775 & vis_psp_o[9]));
assign Snn775 = (~(Non775 & vis_msp_o[9]));
assign Jmn775 = (Uon775 & Bpn775);
assign Bpn775 = (~(Ipn775 & vis_r12_o[11]));
assign Uon775 = (~(Ppn775 & vis_r11_o[11]));
assign Vln775 = (Wpn775 & Dqn775);
assign Dqn775 = (Kqn775 & Rqn775);
assign Rqn775 = (~(Yqn775 & vis_r10_o[11]));
assign Kqn775 = (~(Frn775 & vis_r9_o[11]));
assign Wpn775 = (Nly675 & Mrn775);
assign Mrn775 = (~(Trn775 & vis_r8_o[11]));
assign Pin775 = (~(F2s675 & Vpy675));
assign Vpy675 = (!M2d775);
assign Bin775 = (T3c775 & Asn775);
assign Asn775 = (~(D9k675 & Xxy675));
assign T3c775 = (Cqy675 ^ Hsn775);
assign U4f775 = (~(Osn775 | Moy675));
assign Moy675 = (Ctn775 ? Vsn775 : O1f775);
assign Vsn775 = (Jtn775 & Qtn775);
assign Qtn775 = (Xtn775 & Eun775);
assign Eun775 = (Lun775 & Sun775);
assign Sun775 = (~(Lnn775 & vis_r14_o[8]));
assign Lun775 = (Zun775 & Gvn775);
assign Gvn775 = (~(Gon775 & vis_psp_o[6]));
assign Zun775 = (~(Non775 & vis_msp_o[6]));
assign Xtn775 = (Nvn775 & Uvn775);
assign Uvn775 = (~(Ipn775 & vis_r12_o[8]));
assign Nvn775 = (~(Ppn775 & vis_r11_o[8]));
assign Jtn775 = (Bwn775 & Iwn775);
assign Iwn775 = (Pwn775 & Wwn775);
assign Wwn775 = (~(Yqn775 & vis_r10_o[8]));
assign Pwn775 = (~(Frn775 & vis_r9_o[8]));
assign Bwn775 = (Zdy675 & Dxn775);
assign Dxn775 = (~(Trn775 & vis_r8_o[8]));
assign O1f775 = (!Ewl675);
assign Osn775 = (Wp1l85 ? Rxn775 : Kxn775);
assign Wp1l85 = (~(Yxn775 ^ Kjn775));
assign Yxn775 = (~(Fyn775 & Myn775));
assign Myn775 = (Tyn775 & Azn775);
assign Azn775 = (~(Hzn775 & Fzi675));
assign Tyn775 = (Aln775 | W5f775);
assign Fyn775 = (Ozn775 & Vzn775);
assign Vzn775 = (~(Qgi675 & Fkn775));
assign Ozn775 = (Bx8775 | C0o775);
assign J1n775 = (J0o775 & Q0o775);
assign Q0o775 = (~(X0o775 | Lbe775));
assign Lbe775 = (~(E1o775 | Vwy675));
assign E1o775 = (Qt1l85 ? Rxn775 : Kxn775);
assign Qt1l85 = (~(L1o775 ^ Kjn775));
assign L1o775 = (~(S1o775 & Z1o775));
assign Z1o775 = (~(Pui675 & Fkn775));
assign S1o775 = (G2o775 & Tkn775);
assign G2o775 = (Aln775 | Nce775);
assign X0o775 = (Jhe775 | Qqc775);
assign Qqc775 = (~(N2o775 | Apy675));
assign N2o775 = (Dq1l85 ? Rxn775 : Kxn775);
assign Dq1l85 = (~(U2o775 ^ Kjn775));
assign U2o775 = (~(B3o775 & I3o775));
assign I3o775 = (P3o775 & W3o775);
assign W3o775 = (~(Hzn775 & Xwi675));
assign P3o775 = (Aln775 | Gsc775);
assign B3o775 = (D4o775 & K4o775);
assign K4o775 = (~(Fkn775 & Cei675));
assign D4o775 = (~(Fzi675 & R4o775));
assign Jhe775 = (~(Y4o775 | Cxy675));
assign Cxy675 = (Oln775 ? Dee775 : F5o775);
assign Dee775 = (!U1m675);
assign F5o775 = (M5o775 & T5o775);
assign T5o775 = (A6o775 & H6o775);
assign H6o775 = (O6o775 & V6o775);
assign V6o775 = (~(Lnn775 & vis_r14_o[12]));
assign O6o775 = (C7o775 & J7o775);
assign J7o775 = (~(Gon775 & vis_psp_o[10]));
assign C7o775 = (~(Non775 & vis_msp_o[10]));
assign A6o775 = (Q7o775 & X7o775);
assign X7o775 = (~(Ipn775 & vis_r12_o[12]));
assign Q7o775 = (~(Ppn775 & vis_r11_o[12]));
assign M5o775 = (E8o775 & L8o775);
assign L8o775 = (S8o775 & Z8o775);
assign Z8o775 = (~(Yqn775 & vis_r10_o[12]));
assign S8o775 = (~(Frn775 & vis_r9_o[12]));
assign E8o775 = (Gly675 & G9o775);
assign G9o775 = (~(Trn775 & vis_r8_o[12]));
assign Y4o775 = (Jt1l85 ? Rxn775 : Kxn775);
assign Jt1l85 = (~(N9o775 ^ Kjn775));
assign N9o775 = (~(U9o775 & Bao775));
assign Bao775 = (~(Lti675 & Fkn775));
assign U9o775 = (Iao775 & Tkn775);
assign Iao775 = (Aln775 | Lie775);
assign J0o775 = (Pao775 & Avd775);
assign Avd775 = (Wao775 | Tvy675);
assign Wao775 = (Lu1l85 ? Rxn775 : Kxn775);
assign Lu1l85 = (~(Dbo775 ^ Kjn775));
assign Dbo775 = (~(Kbo775 & Rbo775));
assign Rbo775 = (~(Fzi675 & Fkn775));
assign Kbo775 = (Ybo775 & Tkn775);
assign Ybo775 = (Aln775 | Jwd775);
assign Pao775 = (~(Q9f775 | I6e775));
assign I6e775 = (~(Fco775 | Owy675));
assign Fco775 = (Xt1l85 ? Rxn775 : Kxn775);
assign Xt1l85 = (~(Mco775 ^ Kjn775));
assign Mco775 = (~(Tco775 & Ado775));
assign Ado775 = (~(Tvi675 & Fkn775));
assign Tco775 = (Hdo775 & Tkn775);
assign Hdo775 = (Aln775 | K7e775);
assign Q9f775 = (~(Odo775 | Hwy675));
assign Odo775 = (Su1l85 ? Rxn775 : Kxn775);
assign Su1l85 = (~(Vdo775 ^ Kjn775));
assign Vdo775 = (~(Ceo775 & Jeo775));
assign Jeo775 = (~(Xwi675 & Fkn775));
assign Ceo775 = (Qeo775 & Tkn775);
assign Qeo775 = (Aln775 | Saf775);
assign Ixm775 = (Xeo775 & Efo775);
assign Efo775 = (Lfo775 & Sfo775);
assign Sfo775 = (Zfo775 & Ggo775);
assign Ggo775 = (Ngo775 & Ugo775);
assign Ugo775 = (~(F1e775 | Eqd775));
assign Eqd775 = (~(Bho775 | Mvy675));
assign Bho775 = (Zu1l85 ? Rxn775 : Kxn775);
assign Zu1l85 = (~(Iho775 ^ Kjn775));
assign Iho775 = (~(Pho775 & Who775));
assign Who775 = (~(J0j675 & Fkn775));
assign Pho775 = (Dio775 & Tkn775);
assign Dio775 = (Aln775 | Grd775);
assign F1e775 = (~(Kio775 | Awy675));
assign Awy675 = (Ctn775 ? Rio775 : Zxd775);
assign Rio775 = (Yio775 & Fjo775);
assign Fjo775 = (Mjo775 & Tjo775);
assign Tjo775 = (Ako775 & Hko775);
assign Hko775 = (~(Lnn775 & vis_r14_o[16]));
assign Ako775 = (Oko775 & Vko775);
assign Vko775 = (~(Gon775 & vis_psp_o[14]));
assign Oko775 = (~(Non775 & vis_msp_o[14]));
assign Mjo775 = (Clo775 & Jlo775);
assign Jlo775 = (~(Ipn775 & vis_r12_o[16]));
assign Clo775 = (~(Ppn775 & vis_r11_o[16]));
assign Yio775 = (Qlo775 & Xlo775);
assign Xlo775 = (Emo775 & Lmo775);
assign Lmo775 = (~(Yqn775 & vis_r10_o[16]));
assign Emo775 = (~(Frn775 & vis_r9_o[16]));
assign Qlo775 = (Eky675 & Smo775);
assign Smo775 = (~(Trn775 & vis_r8_o[16]));
assign Zxd775 = (!M7m675);
assign Kio775 = (Eu1l85 ? Rxn775 : Kxn775);
assign Eu1l85 = (~(Zmo775 ^ Kjn775));
assign Zmo775 = (~(Gno775 & Nno775));
assign Nno775 = (~(Byi675 & Fkn775));
assign Gno775 = (Uno775 & Tkn775);
assign Uno775 = (Aln775 | H2e775);
assign H2e775 = (!Boo775);
assign Ngo775 = (~(Qbd775 | Mgd775));
assign Mgd775 = (~(Ioo775 | Ruy675));
assign Ioo775 = (Bw1l85 ? Rxn775 : Kxn775);
assign Bw1l85 = (~(Poo775 ^ Kjn775));
assign Poo775 = (~(Woo775 & Dpo775));
assign Dpo775 = (~(R2j675 & Fkn775));
assign Woo775 = (Kpo775 & Tkn775);
assign Kpo775 = (Aln775 | Ohd775);
assign Ohd775 = (!Rpo775);
assign Qbd775 = (~(Ypo775 | Kuy675));
assign Ypo775 = (Nv1l85 ? Rxn775 : Kxn775);
assign Nv1l85 = (~(Fqo775 ^ Kjn775));
assign Fqo775 = (~(Mqo775 & Tqo775));
assign Tqo775 = (~(V3j675 & Fkn775));
assign Mqo775 = (Aro775 & Tkn775);
assign Aro775 = (Aln775 | Scd775);
assign Scd775 = (!Hro775);
assign Zfo775 = (Oro775 & Uec775);
assign Uec775 = (Vro775 | Bty675);
assign Vro775 = (As1l85 ? Rxn775 : Kxn775);
assign As1l85 = (Rgc775 ? Jso775 : Cso775);
assign Oro775 = (~(Glc775 | Ild775));
assign Ild775 = (~(Qso775 | Fvy675));
assign Qso775 = (Gv1l85 ? Rxn775 : Kxn775);
assign Gv1l85 = (~(Xso775 ^ Kjn775));
assign Xso775 = (~(Eto775 & Lto775));
assign Lto775 = (~(N1j675 & Fkn775));
assign Eto775 = (Sto775 & Tkn775);
assign Sto775 = (Aln775 | Kmd775);
assign Glc775 = (~(Zto775 | Ity675));
assign Ity675 = (Ctn775 ? Guo775 : Mhc775);
assign Guo775 = (Nuo775 & Uuo775);
assign Uuo775 = (Bvo775 & Ivo775);
assign Ivo775 = (Pvo775 & Wvo775);
assign Wvo775 = (~(Lnn775 & vis_r14_o[25]));
assign Pvo775 = (Dwo775 & Kwo775);
assign Kwo775 = (~(Gon775 & vis_psp_o[23]));
assign Dwo775 = (~(Non775 & vis_msp_o[23]));
assign Bvo775 = (Rwo775 & Ywo775);
assign Ywo775 = (~(Ipn775 & vis_r12_o[25]));
assign Rwo775 = (~(Ppn775 & vis_r11_o[25]));
assign Nuo775 = (Fxo775 & Mxo775);
assign Mxo775 = (Txo775 & Ayo775);
assign Ayo775 = (~(Yqn775 & vis_r10_o[25]));
assign Txo775 = (~(Frn775 & vis_r9_o[25]));
assign Fxo775 = (Mhy675 & Hyo775);
assign Hyo775 = (~(Trn775 & vis_r8_o[25]));
assign Mhc775 = (!Hkm675);
assign Zto775 = (Tr1l85 ? Rxn775 : Kxn775);
assign Tr1l85 = (Wmc775 ? Jso775 : Cso775);
assign Lfo775 = (Oyo775 & Vyo775);
assign Vyo775 = (Czo775 & Dab775);
assign Dab775 = (Jzo775 & Qzo775);
assign Qzo775 = (Xzo775 & E0p775);
assign E0p775 = (Cdb775 | L0p775);
assign Xzo775 = (~(Tz1l85[1] | S0p775));
assign S0p775 = (Z0p775 & G1p775);
assign G1p775 = (~(X0a775 | N1p775));
assign Z0p775 = (vis_control_o & U1p775);
assign Jzo775 = (B2p775 & I2p775);
assign I2p775 = (Yuy675 ? W2p775 : P2p775);
assign W2p775 = (~(Ifc775 & Hs1l85));
assign P2p775 = (D3p775 & K3p775);
assign D3p775 = (Hs1l85 ? R3p775 : Ocb775);
assign Hs1l85 = (~(Y3p775 ^ Kjn775));
assign Y3p775 = (~(F4p775 & M4p775));
assign M4p775 = (~(Lti675 & T4p775));
assign F4p775 = (A5p775 & H5p775);
assign H5p775 = (Aln775 | L0p775);
assign A5p775 = (~(T7i675 & Fkn775));
assign B2p775 = (O5p775 & V5p775);
assign V5p775 = (~(Mbb775 & Sy1l85[1]));
assign O5p775 = (~(C6p775 & vis_ipsr_o[1]));
assign Czo775 = (~(J6p775 | N6d775));
assign N6d775 = (~(Q6p775 | Duy675));
assign Q6p775 = (Uv1l85 ? Rxn775 : Kxn775);
assign Uv1l85 = (~(X6p775 ^ Kjn775));
assign X6p775 = (~(E7p775 & L7p775));
assign L7p775 = (Tli675 ? Z7p775 : S7p775);
assign S7p775 = (~(Fkn775 & Fd9775));
assign E7p775 = (G8p775 & Tkn775);
assign G8p775 = (Aln775 | P7d775);
assign J6p775 = (N8p775 & U8p775);
assign U8p775 = (~(B9p775 & I9p775));
assign I9p775 = (P9p775 & W9p775);
assign W9p775 = (Dap775 & Kap775);
assign Kap775 = (Rap775 & Kmd775);
assign Rap775 = (~(Rpo775 | Hro775));
assign Dap775 = (~(Yap775 | Fbp775));
assign P9p775 = (Mbp775 & Tbp775);
assign Tbp775 = (Acp775 & Rgc775);
assign Acp775 = (~(Hcp775 | Ocp775));
assign Mbp775 = (~(Vcp775 | Cdp775));
assign B9p775 = (Jdp775 & Qdp775);
assign Qdp775 = (Xdp775 & Eep775);
assign Eep775 = (Lep775 & Saf775);
assign Lep775 = (~(Boo775 | Sep775));
assign Xdp775 = (~(Zep775 | Gfp775));
assign Jdp775 = (Nfp775 & Ufp775);
assign Ufp775 = (~(Bgp775 | Igp775));
assign Nfp775 = (~(Pgp775 | Wgp775));
assign Oyo775 = (Dhp775 & G0c775);
assign G0c775 = (Khp775 & Rhp775);
assign Rhp775 = (Yhp775 & Fip775);
assign Fip775 = (~(Mbb775 & Sy1l85[7]));
assign Yhp775 = (~(Tz1l85[7] | Gec775));
assign Khp775 = (Mip775 & Tip775);
assign Tip775 = (~(N8p775 & Ajp775));
assign Mip775 = (Toy675 ? Ojp775 : Hjp775);
assign Ojp775 = (~(Ifc775 & Ip1l85));
assign Hjp775 = (Ip1l85 ? Rxn775 : Kxn775);
assign Ip1l85 = (~(Vjp775 ^ Kjn775));
assign Vjp775 = (~(Ckp775 & Jkp775));
assign Jkp775 = (Qkp775 & Xkp775);
assign Xkp775 = (~(Hzn775 & Byi675));
assign Qkp775 = (Aln775 | Elp775);
assign Ckp775 = (Llp775 & Slp775);
assign Slp775 = (~(Fkn775 & Jfi675));
assign Llp775 = (~(J0j675 & R4o775));
assign Dhp775 = (I1c775 & U0c775);
assign U0c775 = (Zlp775 & Gmp775);
assign Gmp775 = (Nmp775 & Ump775);
assign Ump775 = (~(Bnp775 & vis_apsr_o[0]));
assign Nmp775 = (~(Tz1l85[28] | Gec775));
assign Zlp775 = (Inp775 & Pnp775);
assign Pnp775 = (Nsy675 ? Dop775 : Wnp775);
assign Dop775 = (~(Ifc775 & Rq1l85));
assign Wnp775 = (Kop775 & K3p775);
assign Kop775 = (Rq1l85 ? R3p775 : Ocb775);
assign Rq1l85 = (Dz0775 ? Jso775 : Cso775);
assign Inp775 = (Rop775 & Yop775);
assign Yop775 = (Cdb775 | Dz0775);
assign Rop775 = (~(Mbb775 & Sy1l85[28]));
assign I1c775 = (Fpp775 & Mpp775);
assign Mpp775 = (Tpp775 & Aqp775);
assign Aqp775 = (~(N8p775 & Pig775));
assign Tpp775 = (~(Tz1l85[31] | Gec775));
assign Fpp775 = (Hqp775 & Oqp775);
assign Oqp775 = (V2l775 ? Crp775 : Vqp775);
assign Crp775 = (~(Ifc775 & Kq1l85));
assign Vqp775 = (Kq1l85 ? Rxn775 : Kxn775);
assign Kq1l85 = (Pig775 ? Cso775 : Jso775);
assign Hqp775 = (Jrp775 & Qrp775);
assign Qrp775 = (~(vis_apsr_o[3] & Bnp775));
assign Jrp775 = (~(Mbb775 & Sy1l85[31]));
assign Xeo775 = (Xrp775 & Esp775);
assign Esp775 = (Lsp775 & Ssp775);
assign Ssp775 = (Zsp775 & A3d775);
assign A3d775 = (Gtp775 & Ntp775);
assign Ntp775 = (~(C6p775 & vis_ipsr_o[3]));
assign Gtp775 = (~(Tz1l85[3] | Utp775));
assign Utp775 = (Bup775 & M2d775);
assign M2d775 = (Ctn775 ? Iup775 : Gpl675);
assign Iup775 = (~(Pup775 & Wup775));
assign Wup775 = (Dvp775 & Kvp775);
assign Kvp775 = (Rvp775 & Yvp775);
assign Yvp775 = (~(Lnn775 & vis_r14_o[3]));
assign Rvp775 = (Fwp775 & Mwp775);
assign Mwp775 = (~(Gon775 & vis_psp_o[1]));
assign Fwp775 = (~(Non775 & vis_msp_o[1]));
assign Dvp775 = (Twp775 & Axp775);
assign Axp775 = (~(Ipn775 & vis_r12_o[3]));
assign Twp775 = (~(Ppn775 & vis_r11_o[3]));
assign Pup775 = (Hxp775 & Oxp775);
assign Oxp775 = (Vxp775 & Cyp775);
assign Cyp775 = (~(Yqn775 & vis_r10_o[3]));
assign Vxp775 = (~(Frn775 & vis_r9_o[3]));
assign Hxp775 = (Ify675 & Jyp775);
assign Jyp775 = (~(Trn775 & vis_r8_o[3]));
assign Bup775 = (F2s675 ? E9n775 : X8n775);
assign F2s675 = (~(Qyp775 ^ Kjn775));
assign Qyp775 = (~(Xyp775 & Ezp775));
assign Ezp775 = (Lzp775 & Szp775);
assign Szp775 = (So1775 | Zzp775);
assign So1775 = (!Lti675);
assign Lzp775 = (Aln775 | K1d775);
assign Xyp775 = (G0q775 & N0q775);
assign N0q775 = (~(Hai675 & Fkn775));
assign G0q775 = (~(Tvi675 & R4o775));
assign Zsp775 = (O4c775 & Qdb775);
assign Qdb775 = (U0q775 & B1q775);
assign B1q775 = (I1q775 & P1q775);
assign P1q775 = (~(W1q775 & D2q775));
assign D2q775 = (~(N1p775 | Pui675));
assign W1q775 = (U1p775 & vis_primask_o);
assign I1q775 = (~(Tz1l85[0] | Gec775));
assign U0q775 = (K2q775 & R2q775);
assign R2q775 = (~(Y2q775 & Vcb775));
assign Y2q775 = (D9k675 ? E9n775 : X8n775);
assign D9k675 = (~(F3q775 ^ Kjn775));
assign F3q775 = (~(M3q775 & T3q775));
assign T3q775 = (Aln775 | Jdb775);
assign M3q775 = (~(Hsi675 & T4p775));
assign E9n775 = (!Rxn775);
assign X8n775 = (!Kxn775);
assign K2q775 = (~(C6p775 & vis_ipsr_o[0]));
assign O4c775 = (A4q775 & H4q775);
assign H4q775 = (~(vis_apsr_o[2] & Bnp775));
assign A4q775 = (~(Tz1l85[30] | O4q775));
assign O4q775 = (Cqy675 & V4q775);
assign V4q775 = (~(K3p775 & C5q775));
assign C5q775 = (Hsn775 | R3p775);
assign Hsn775 = (!Nak675);
assign Nak675 = (~(J5q775 & Q5q775));
assign J5q775 = (Ocp775 ? E6q775 : X5q775);
assign Lsp775 = (L6q775 & Ruc775);
assign Ruc775 = (S6q775 & Z6q775);
assign Z6q775 = (G7q775 & N7q775);
assign N7q775 = (~(N8p775 & U7q775));
assign G7q775 = (~(Tz1l85[5] | Gec775));
assign S6q775 = (B8q775 & I8q775);
assign I8q775 = (Hpy675 ? W8q775 : P8q775);
assign W8q775 = (~(Ifc775 & No1l85));
assign P8q775 = (D9q775 & K3p775);
assign D9q775 = (No1l85 ? R3p775 : Ocb775);
assign No1l85 = (~(K9q775 ^ Kjn775));
assign K9q775 = (~(R9q775 & Y9q775));
assign Y9q775 = (Faq775 & Maq775);
assign Maq775 = (Gga775 | Zzp775);
assign Gga775 = (!Tvi675);
assign Faq775 = (~(Taq775 & U7q775));
assign R9q775 = (Abq775 & Hbq775);
assign Hbq775 = (~(Fkn775 & Vci675));
assign Abq775 = (~(Byi675 & R4o775));
assign B8q775 = (Obq775 & Vbq775);
assign Vbq775 = (~(Mbb775 & Sy1l85[5]));
assign Obq775 = (~(C6p775 & vis_ipsr_o[5]));
assign L6q775 = (Cxc775 & Gxe775);
assign Gxe775 = (Ccq775 & Jcq775);
assign Jcq775 = (Qcq775 & Xcq775);
assign Xcq775 = (~(Tz1l85[2] | Edq775));
assign Edq775 = (Ldq775 & Sdq775);
assign Sdq775 = (Gvo675 & W1p675);
assign Ldq775 = (N6i675 & V7g775);
assign Qcq775 = (Zdq775 & Geq775);
assign Geq775 = (~(Gec775 & vis_control_o));
assign Zdq775 = (Cdb775 | Neq775);
assign Ccq775 = (Ueq775 & Bfq775);
assign Bfq775 = (Xqy675 ? Pfq775 : Ifq775);
assign Xqy675 = (Oln775 ? Wnl675 : Wfq775);
assign Wfq775 = (~(Dgq775 & Kgq775));
assign Kgq775 = (Rgq775 & Ygq775);
assign Ygq775 = (Fhq775 & Mhq775);
assign Mhq775 = (~(Lnn775 & vis_r14_o[2]));
assign Fhq775 = (Thq775 & Aiq775);
assign Aiq775 = (~(Gon775 & vis_psp_o[0]));
assign Thq775 = (~(Non775 & vis_msp_o[0]));
assign Rgq775 = (Hiq775 & Oiq775);
assign Oiq775 = (~(Ipn775 & vis_r12_o[2]));
assign Hiq775 = (~(Ppn775 & vis_r11_o[2]));
assign Dgq775 = (Viq775 & Cjq775);
assign Cjq775 = (Jjq775 & Qjq775);
assign Qjq775 = (~(Yqn775 & vis_r10_o[2]));
assign Jjq775 = (~(Frn775 & vis_r9_o[2]));
assign Viq775 = (Dgy675 & Xjq775);
assign Xjq775 = (~(Trn775 & vis_r8_o[2]));
assign Pfq775 = (Ekq775 & K3p775);
assign Ekq775 = (Bp1l85 ? R3p775 : Ocb775);
assign Ifq775 = (Ocb775 | Lkq775);
assign Lkq775 = (!Bp1l85);
assign Bp1l85 = (~(Skq775 ^ Kjn775));
assign Skq775 = (~(Zkq775 & Glq775));
assign Glq775 = (Nlq775 & Ulq775);
assign Ulq775 = (Xo0775 | Zzp775);
assign Nlq775 = (Aln775 | Neq775);
assign Zkq775 = (Bmq775 & Imq775);
assign Imq775 = (~(A9i675 & Fkn775));
assign Bmq775 = (~(Pui675 & T4p775));
assign T4p775 = (R4o775 | Pmq775);
assign Pmq775 = (Wmq775 & Dnq775);
assign Dnq775 = (~(Nvg775 | K1z675));
assign Wmq775 = (Sa1775 & Gvo675);
assign Ueq775 = (Knq775 & Rnq775);
assign Rnq775 = (~(Mbb775 & Sy1l85[2]));
assign Knq775 = (~(C6p775 & vis_ipsr_o[2]));
assign Cxc775 = (Ynq775 & Foq775);
assign Foq775 = (Moq775 & Toq775);
assign Toq775 = (~(N8p775 & Apq775));
assign Moq775 = (~(Tz1l85[4] | Gec775));
assign Ynq775 = (Hpq775 & Opq775);
assign Opq775 = (Opy675 ? Cqq775 : Vpq775);
assign Cqq775 = (~(Ifc775 & Uo1l85));
assign Vpq775 = (Jqq775 & K3p775);
assign Jqq775 = (Uo1l85 ? R3p775 : Ocb775);
assign Uo1l85 = (~(Qqq775 ^ Kjn775));
assign Qqq775 = (~(Xqq775 & Erq775));
assign Erq775 = (Lrq775 & Srq775);
assign Srq775 = (X0a775 | Zzp775);
assign Zzp775 = (~(Hzn775 | Zrq775));
assign Zrq775 = (Gvo675 & Gsq775);
assign Gsq775 = (~(Nsq775 & Usq775));
assign Usq775 = (Btq775 & Itq775);
assign Itq775 = (~(Ptq775 & O4p675));
assign Ptq775 = (Wtq775 & Cm2775);
assign Wtq775 = (~(Duq775 & Kuq775));
assign Kuq775 = (Ryf775 | Xza775);
assign Btq775 = (~(Mwo675 & Vs9775));
assign Vs9775 = (Zx6775 | Sh1775);
assign Nsq775 = (Ruq775 & Yuq775);
assign Yuq775 = (~(Fvq775 & Ub1775));
assign Ruq775 = (Yyf775 | Cg8775);
assign Lrq775 = (~(Taq775 & Apq775));
assign Xqq775 = (Mvq775 & Tvq775);
assign Tvq775 = (~(Obi675 & Fkn775));
assign Mvq775 = (~(Xwi675 & R4o775));
assign R4o775 = (~(C0o775 & Awq775));
assign Awq775 = (~(Gvo675 & Hwq775));
assign Hwq775 = (~(Owq775 & Vwq775));
assign Vwq775 = (~(Cxq775 & Cg8775));
assign Cxq775 = (~(Jxq775 & Qxq775));
assign Qxq775 = (~(Xxq775 & Xza775));
assign Owq775 = (Eyq775 & Lyq775);
assign Lyq775 = (~(Kny675 & Syq775));
assign Syq775 = (~(O2l775 & Zyq775));
assign Zyq775 = (Zry675 | F3p675);
assign Eyq775 = (~(Bvh675 & Gzq775));
assign Gzq775 = (~(Wdl775 & Nzq775));
assign Nzq775 = (~(Fvq775 & Mwo675));
assign Hpq775 = (Uzq775 & B0r775);
assign B0r775 = (~(Mbb775 & Sy1l85[4]));
assign Uzq775 = (~(C6p775 & vis_ipsr_o[4]));
assign C6p775 = (I0r775 & U1p775);
assign I0r775 = (~(Xo0775 | Xwi675));
assign Xo0775 = (!Hsi675);
assign Xrp775 = (P0r775 & W0r775);
assign W0r775 = (D1r775 & D9c775);
assign D9c775 = (K1r775 & R1r775);
assign R1r775 = (Y1r775 & F2r775);
assign F2r775 = (~(Bnp775 & vis_apsr_o[1]));
assign Bnp775 = (Wig775 & U1p775);
assign U1p775 = (M2r775 & Ssb775);
assign M2r775 = (Gvo675 & T2r775);
assign Wig775 = (~(Pui675 | Xwi675));
assign Y1r775 = (~(Tz1l85[29] | Gec775));
assign K1r775 = (A3r775 & H3r775);
assign H3r775 = (Gsy675 ? V3r775 : O3r775);
assign V3r775 = (~(Ifc775 & Yq1l85));
assign O3r775 = (C4r775 & K3p775);
assign C4r775 = (Yq1l85 ? R3p775 : Ocb775);
assign Yq1l85 = (Ft0775 ? Cso775 : Jso775);
assign A3r775 = (J4r775 & Q4r775);
assign Q4r775 = (~(N8p775 & Ft0775));
assign J4r775 = (~(Mbb775 & Sy1l85[29]));
assign D1r775 = (~(Hbc775 | T0f775));
assign T0f775 = (~(X4r775 & E5r775));
assign E5r775 = (L5r775 & S5r775);
assign S5r775 = (~(N8p775 & Z5r775));
assign L5r775 = (~(Tz1l85[9] | Gec775));
assign X4r775 = (G6r775 & N6r775);
assign N6r775 = (~(Mbb775 & Sy1l85[9]));
assign G6r775 = (Yny675 ? B7r775 : U6r775);
assign Yny675 = (Ctn775 ? I7r775 : F0f775);
assign I7r775 = (P7r775 & W7r775);
assign W7r775 = (D8r775 & K8r775);
assign K8r775 = (R8r775 & Y8r775);
assign Y8r775 = (~(Lnn775 & vis_r14_o[9]));
assign R8r775 = (F9r775 & M9r775);
assign M9r775 = (~(Gon775 & vis_psp_o[7]));
assign F9r775 = (~(Non775 & vis_msp_o[7]));
assign D8r775 = (T9r775 & Aar775);
assign Aar775 = (~(Ipn775 & vis_r12_o[9]));
assign T9r775 = (~(Ppn775 & vis_r11_o[9]));
assign P7r775 = (Har775 & Oar775);
assign Oar775 = (Var775 & Cbr775);
assign Cbr775 = (~(Yqn775 & vis_r10_o[9]));
assign Var775 = (~(Frn775 & vis_r9_o[9]));
assign Har775 = (Sdy675 & Jbr775);
assign Jbr775 = (~(Trn775 & vis_r8_o[9]));
assign F0f775 = (!Oxl675);
assign B7r775 = (~(Ifc775 & Pp1l85));
assign U6r775 = (Qbr775 & K3p775);
assign Qbr775 = (Pp1l85 ? R3p775 : Ocb775);
assign Pp1l85 = (~(Xbr775 ^ Kjn775));
assign Xbr775 = (~(Ecr775 & Lcr775));
assign Lcr775 = (Scr775 & Zcr775);
assign Zcr775 = (~(Hzn775 & J0j675));
assign Hzn775 = (Gvo675 & Gdr775);
assign Gdr775 = (~(Ndr775 & Udr775));
assign Udr775 = (Ezo675 ? Ier775 : Ber775);
assign Ier775 = (~(Per775 & A3z675));
assign Ber775 = (Pyl775 | Xuf775);
assign Ndr775 = (Wer775 & Dfr775);
assign Dfr775 = (~(Kfr775 & Ssb775));
assign Ssb775 = (~(Bbg775 | Bvh675));
assign Kfr775 = (Rcg775 & Kny675);
assign Wer775 = (~(Rfr775 & Yfr775));
assign Yfr775 = (Fgr775 | Per775);
assign Fgr775 = (Zrj775 | Ezo675);
assign Scr775 = (~(Taq775 & Z5r775));
assign Ecr775 = (Mgr775 & Tgr775);
assign Tgr775 = (~(Xhi675 & Fkn775));
assign Mgr775 = (B49775 | C0o775);
assign Hbc775 = (~(Ahr775 & Hhr775));
assign Hhr775 = (Ohr775 & Vhr775);
assign Vhr775 = (~(N8p775 & Cir775));
assign Ohr775 = (~(Tz1l85[27] | Gec775));
assign Ahr775 = (Jir775 & Qir775);
assign Qir775 = (~(Mbb775 & Sy1l85[27]));
assign Jir775 = (Usy675 ? Ejr775 : Xir775);
assign Ejr775 = (~(Ifc775 & Fr1l85));
assign Xir775 = (Ljr775 & K3p775);
assign Ljr775 = (Fr1l85 ? R3p775 : Ocb775);
assign Fr1l85 = (Cir775 ? Cso775 : Jso775);
assign P0r775 = (Sjr775 & Xfg775);
assign Xfg775 = (Zjr775 & Gkr775);
assign Gkr775 = (Nkr775 & Ukr775);
assign Ukr775 = (~(Mbb775 & Sy1l85[23]));
assign Nkr775 = (~(Tz1l85[23] | Gec775));
assign Zjr775 = (Blr775 & Ilr775);
assign Ilr775 = (Cdb775 | Plr775);
assign Blr775 = (Wty675 ? Dmr775 : Wlr775);
assign Dmr775 = (~(Ifc775 & Os1l85));
assign Wlr775 = (Os1l85 ? Rxn775 : Kxn775);
assign Os1l85 = (~(Kmr775 ^ Kjn775));
assign Kmr775 = (Rmr775 | Ymr775);
assign Ymr775 = (Joi675 ? Mnr775 : Fnr775);
assign Fnr775 = (Fkn775 & Fd9775);
assign Rmr775 = (~(Tnr775 & Tkn775));
assign Tnr775 = (Aln775 | Plr775);
assign Sjr775 = (Dse775 & Knc775);
assign Knc775 = (Aor775 & Hor775);
assign Hor775 = (Oor775 & Vor775);
assign Vor775 = (~(Mbb775 & Sy1l85[24]));
assign Oor775 = (~(Tz1l85[24] | Gec775));
assign Aor775 = (Cpr775 & Jpr775);
assign Jpr775 = (~(N8p775 & Qpr775));
assign Cpr775 = (Pty675 ? Eqr775 : Xpr775);
assign Eqr775 = (~(Ifc775 & Mr1l85));
assign Xpr775 = (Mr1l85 ? Rxn775 : Kxn775);
assign Mr1l85 = (Qpr775 ? Cso775 : Jso775);
assign Cso775 = (~(Q5q775 & E6q775));
assign E6q775 = (~(Taq775 & Kjn775));
assign Jso775 = (~(Q5q775 & X5q775));
assign Q5q775 = (Lqr775 & Sqr775);
assign Sqr775 = (X5q775 | Taq775);
assign Taq775 = (!Aln775);
assign X5q775 = (Zqr775 | Kjn775);
assign Lqr775 = (~(Kjn775 & Zqr775));
assign Zqr775 = (~(Z7p775 & Tkn775));
assign Tkn775 = (Fd9775 | C0o775);
assign Z7p775 = (!Mnr775);
assign Mnr775 = (Fkn775 & A5j675);
assign Dse775 = (Grr775 & Nrr775);
assign Nrr775 = (Urr775 & Bsr775);
assign Bsr775 = (~(Mbb775 & Sy1l85[10]));
assign Mbb775 = (Gvo675 & Isr775);
assign Isr775 = (Psr775 | Gvg775);
assign Psr775 = (N0p675 ? Ex6775 : Wsr775);
assign Wsr775 = (~(Dtr775 & Ktr775));
assign Ktr775 = (Wbg775 | Rto675);
assign Dtr775 = (~(Rtr775 | Ytr775));
assign Urr775 = (~(Tz1l85[10] | Gec775));
assign Gec775 = (!M3c775);
assign M3c775 = (~(Fur775 & Gvo675));
assign Fur775 = (Dny675 & Rto675);
assign Grr775 = (Mur775 & Tur775);
assign Tur775 = (Cdb775 | Avr775);
assign Cdb775 = (!N8p775);
assign N8p775 = (Gvo675 & Hvr775);
assign Hvr775 = (~(Ovr775 & Tsf775));
assign Ovr775 = (~(Psk775 & Vvr775));
assign Mur775 = (Qxy675 ? Jwr775 : Cwr775);
assign Jwr775 = (~(Ifc775 & Vs1l85));
assign Ifc775 = (!Ocb775);
assign Cwr775 = (Vs1l85 ? Rxn775 : Kxn775);
assign Vs1l85 = (~(Qwr775 ^ Kjn775));
assign Kjn775 = (~(Gvo675 & Xwr775));
assign Xwr775 = (~(Exr775 & Lxr775));
assign Lxr775 = (Sxr775 & Zxr775);
assign Zxr775 = (~(Gyr775 & Xza775));
assign Gyr775 = (~(Nyr775 & Uyr775));
assign Uyr775 = (~(Bzr775 & Vxo675));
assign Sxr775 = (Izr775 & X4z675);
assign X4z675 = (~(Pzr775 & Wzr775));
assign Izr775 = (~(D0s775 & Ytr775));
assign D0s775 = (~(Jbk775 | Cm2775));
assign Exr775 = (J4z675 & K0s775);
assign K0s775 = (~(Bzr775 & Uag775));
assign J4z675 = (R0s775 & Y0s775);
assign Y0s775 = (Wxf775 | Eta775);
assign R0s775 = (F1s775 & M1s775);
assign M1s775 = (O2l775 | Cm2775);
assign O2l775 = (!T1s775);
assign F1s775 = (~(M6g775 & Kny675));
assign Qwr775 = (~(A2s775 & H2s775));
assign H2s775 = (Amf775 | C0o775);
assign C0o775 = (~(O2s775 & Gvo675));
assign O2s775 = (~(Oya775 | Rxg775));
assign A2s775 = (V2s775 & C3s775);
assign C3s775 = (Aln775 | Avr775);
assign Aln775 = (~(Gvo675 & J3s775));
assign J3s775 = (~(Q3s775 & X3s775));
assign X3s775 = (E4s775 & L4s775);
assign L4s775 = (~(S4s775 & Uag775));
assign S4s775 = (Pxf775 & Ezo675);
assign E4s775 = (~(Z4s775 | Bzr775));
assign Q3s775 = (G5s775 & N5s775);
assign N5s775 = (Yyf775 | Rxg775);
assign G5s775 = (U5s775 & B6s775);
assign B6s775 = (~(I6s775 & Lx6775));
assign I6s775 = (~(Xuf775 | Del775));
assign U5s775 = (~(Rto675 & P6s775));
assign P6s775 = (~(W6s775 & D7s775));
assign D7s775 = (K7s775 | I6l775);
assign W6s775 = (R7s775 & Pyl775);
assign R7s775 = (~(Ezo675 & Y7s775));
assign Y7s775 = (U50775 | N0p675);
assign V2s775 = (~(Eji675 & Fkn775));
assign Fkn775 = (F8s775 & M8s775);
assign M8s775 = (Kny675 & Y1z675);
assign F8s775 = (Gvo675 & N0p675);
assign Rxn775 = (R3p775 & K3p775);
assign R3p775 = (T8s775 & A9s775);
assign A9s775 = (~(H9s775 & Rto675));
assign H9s775 = (O9s775 & K1z675);
assign O9s775 = (D1z675 | O0g775);
assign T8s775 = (Pyl775 | I6l775);
assign Pyl775 = (!O0g775);
assign Kxn775 = (K3p775 & Ocb775);
assign Ocb775 = (~(V9s775 & Bzr775));
assign Bzr775 = (N0p675 & D1z675);
assign V9s775 = (Gvo675 & V0g775);
assign K3p775 = (~(Gvo675 & Cas775));
assign Cas775 = (~(Jas775 & Qas775));
assign Qas775 = (Xas775 & Kp3775);
assign Jas775 = (Ebs775 & Lbs775);
assign Lbs775 = (~(Eck775 & Lrh675));
assign Ebs775 = (F3p675 ? Zbs775 : Sbs775);
assign Zbs775 = (Q6b775 | Pw9775);
assign Sbs775 = (Veg775 | N0p675);
assign Ovk775 = (~(Gcs775 & Ncs775));
assign Gcs775 = (Ucs775 & M53775);
assign Ucs775 = (Dqg775 | Bds775);
assign Bds775 = (Ids775 & Pds775);
assign Ids775 = (~(Ty2775 | Tli675));
assign Avk775 = (Wds775 & Des775);
assign Des775 = (~(Kes775 & Wk0775));
assign Kes775 = (~(Yyf775 | K1z675));
assign Wds775 = (~(Res775 & Hph675));
assign Res775 = (~(Ep0775 | O4p675));
assign Muk775 = (Yes775 & Ffs775);
assign Ffs775 = (M2k775 | Rto675);
assign Yes775 = (Mfs775 & Tfs775);
assign Tfs775 = (~(Vwj775 & Ags775));
assign Ags775 = (~(Hgs775 & Lki675));
assign Hgs775 = (M53775 ? Ogs775 : Eji675);
assign Mfs775 = (~(Vgs775 & Chs775));
assign Ytk775 = (Jhs775 & Qhs775);
assign Qhs775 = (Xhs775 & Eis775);
assign Eis775 = (~(Xxq775 & Lis775));
assign Xhs775 = (Sis775 & Zis775);
assign Zis775 = (~(Gjs775 & Njs775));
assign Njs775 = (~(Ujs775 & Bks775));
assign Bks775 = (Iks775 & Pks775);
assign Pks775 = (R1z675 | U50775);
assign Iks775 = (Wks775 | F3p675);
assign Ujs775 = (Mwo675 & Dls775);
assign Dls775 = (Y1z675 | N0p675);
assign Sis775 = (~(Kls775 & Rls775));
assign Rls775 = (~(Yls775 & Fms775));
assign Fms775 = (Mms775 & Tms775);
assign Tms775 = (~(Ans775 & Hns775));
assign Ans775 = (~(V8p675 | Rto675));
assign Mms775 = (~(Ons775 & Vns775));
assign Vns775 = (~(W1p675 & Cos775));
assign Cos775 = (~(Jos775 & Qos775));
assign Yls775 = (Xos775 & Eps775);
assign Eps775 = (~(A3k775 & Zx6775));
assign Xos775 = (~(Lps775 & Q91775));
assign Jhs775 = (Sps775 & Zps775);
assign Sps775 = (Gqs775 & Nqs775);
assign Nqs775 = (~(Vjb775 & Yuj775));
assign Gqs775 = (C8g775 | Fkg775);
assign D1s675 = (Uqs775 & Brs775);
assign Brs775 = (~(Irs775 & Prs775));
assign Prs775 = (Wrs775 & Dss775);
assign Dss775 = (Kss775 & Rss775);
assign Rss775 = (Yss775 & Iw9775);
assign Yss775 = (~(Fts775 & Rvb775));
assign Kss775 = (Mts775 & Tts775);
assign Tts775 = (~(Aus775 & Hus775));
assign Hus775 = (Zqi675 | Ous775);
assign Mts775 = (~(Vus775 & U50775));
assign Vus775 = (My9775 | Osg775);
assign Wrs775 = (Cvs775 & Jvs775);
assign Jvs775 = (Qvs775 & Xvs775);
assign Xvs775 = (~(Ews775 & Y1z675));
assign Ews775 = (Jf9775 | Eck775);
assign Qvs775 = (Lws775 | Tc3775);
assign Cvs775 = (Sws775 & Zws775);
assign Zws775 = (~(Gxs775 & Bek775));
assign Sws775 = (~(Nxs775 & Uxs775));
assign Uxs775 = (~(Bys775 & Iys775));
assign Iys775 = (Pys775 & Wys775);
assign Wys775 = (~(Rpi675 | Qgi675));
assign Pys775 = (~(Dzs775 | Kzs775));
assign Dzs775 = (~(Tc3775 | Qpk775));
assign Qpk775 = (Rzs775 & Yzs775);
assign Rzs775 = (~(Vci675 | Jfi675));
assign Bys775 = (F0t775 & Izk775);
assign F0t775 = (~(Ye0775 | Ty2775));
assign Irs775 = (M0t775 & T0t775);
assign T0t775 = (A1t775 & H1t775);
assign H1t775 = (O1t775 & V1t775);
assign V1t775 = (~(Rpi675 & C2t775));
assign C2t775 = (~(J2t775 & Q2t775));
assign Q2t775 = (X2t775 & E3t775);
assign E3t775 = (~(Aus775 & L3t775));
assign L3t775 = (~(S3t775 & Z3t775));
assign Z3t775 = (G4t775 & Tc3775);
assign G4t775 = (~(N4t775 & Kzs775));
assign N4t775 = (~(A9l775 | Qgi675));
assign S3t775 = (U4t775 & B5t775);
assign B5t775 = (~(Xhi675 & I5t775));
assign I5t775 = (~(P5t775 & W5t775));
assign W5t775 = (Lyj775 | Eji675);
assign X2t775 = (~(D6t775 & Bvh675));
assign J2t775 = (K6t775 & R6t775);
assign R6t775 = (A9l775 | J6b775);
assign K6t775 = (~(Izk775 & N9a775));
assign O1t775 = (~(Uo9775 & Xhi675));
assign A1t775 = (Y6t775 & F7t775);
assign F7t775 = (~(Os9775 & T2r775));
assign Y6t775 = (~(Eck775 & M7t775));
assign M0t775 = (T7t775 & A8t775);
assign A8t775 = (~(H8t775 | O8t775));
assign O8t775 = (Zck775 & Srj775);
assign T7t775 = (~(V8t775 | C9t775));
assign C9t775 = (F3p675 ? J9t775 : Z8a775);
assign J9t775 = (~(Q6b775 | Ibg775));
assign V8t775 = (O4p675 ? Q9t775 : Osg775);
assign Q9t775 = (~(X9t775 & Eat775));
assign Eat775 = (Lat775 & Sat775);
assign Sat775 = (~(Zat775 & My9775));
assign Zat775 = (~(O6a775 | Kls775));
assign Lat775 = (~(Eh1775 & Iso675));
assign X9t775 = (Gbt775 & Nbt775);
assign Nbt775 = (~(Frg775 & F6g775));
assign Gbt775 = (Ryf775 | Bvh675);
assign Uqs775 = (O4p675 | hready_i);
assign W0s675 = (Bct775 ? Iw1l85[3] : Ubt775);
assign Ubt775 = (~(Ict775 & Pct775));
assign Pct775 = (~(Qgi675 & Wct775));
assign Wct775 = (Ddt775 | Kdt775);
assign Kdt775 = (Rdt775 & Lki675);
assign P0s675 = (~(Ydt775 & Fet775));
assign Fet775 = (Met775 & Tet775);
assign Tet775 = (~(Aft775 & Sy1l85[30]));
assign Met775 = (Hft775 & Oft775);
assign Hft775 = (Vft775 | H4c775);
assign H4c775 = (Cgt775 & Jgt775);
assign Jgt775 = (Qgt775 & Xgt775);
assign Xgt775 = (~(Eht775 & Lht775));
assign Qgt775 = (Sht775 & Zht775);
assign Sht775 = (Git775 | Nit775);
assign Cgt775 = (Uit775 & Bjt775);
assign Bjt775 = (~(Ijt775 & Pjt775));
assign Uit775 = (~(Wjt775 & Dkt775));
assign Ydt775 = (Kkt775 & Rkt775);
assign Rkt775 = (~(E52l85[29] & Ykt775));
assign Kkt775 = (~(vis_pc_o[29] & P60775));
assign I0s675 = (Flt775 | Mlt775);
assign Mlt775 = (~(Olg775 | F3p675));
assign Flt775 = (hready_i ? Tlt775 : Vxo675);
assign Tlt775 = (~(Amt775 & Hmt775));
assign Hmt775 = (Omt775 & Vmt775);
assign Vmt775 = (Cnt775 & Jnt775);
assign Jnt775 = (~(Qnt775 & Xnt775));
assign Xnt775 = (!Eot775);
assign Cnt775 = (~(Lot775 & Y1z675));
assign Lot775 = (~(Sot775 & Zot775));
assign Zot775 = (~(Gpt775 & Gjs775));
assign Gpt775 = (~(Yyf775 | W1p675));
assign Omt775 = (Npt775 & Upt775);
assign Upt775 = (~(Bqt775 & M71775));
assign Bqt775 = (~(Iqt775 & Pqt775));
assign Pqt775 = (Ky8775 | Tc3775);
assign Iqt775 = (Wqt775 & Drt775);
assign Drt775 = (~(D6t775 & Q89775));
assign Wqt775 = (~(Hns775 & A3z675));
assign Hns775 = (Krt775 & Vsg775);
assign Krt775 = (~(Te1775 | Q91775));
assign Npt775 = (~(Rrt775 & E5z675));
assign Rrt775 = (~(Yrt775 & Fst775));
assign Fst775 = (Mst775 & Pub775);
assign Mst775 = (Tst775 & Att775);
assign Yrt775 = (Htt775 & Ott775);
assign Ott775 = (~(Vtt775 & Cut775));
assign Htt775 = (Jut775 & Rny675);
assign Jut775 = (~(Rvb775 & Qut775));
assign Qut775 = (Mdg775 | Xut775);
assign Amt775 = (Evt775 & Lvt775);
assign Lvt775 = (Svt775 & Zvt775);
assign Zvt775 = (~(Wc1775 & Gwt775));
assign Gwt775 = (~(Nwt775 & Uwt775));
assign Uwt775 = (Bxt775 & Ixt775);
assign Ixt775 = (~(Tli675 & Pxt775));
assign Pxt775 = (Wxt775 | Dyt775);
assign Dyt775 = (Lki675 ? Kyt775 : Nxs775);
assign Kyt775 = (~(Ryt775 | Cm2775));
assign Wxt775 = (~(Yyt775 & Fzt775));
assign Fzt775 = (~(Mzt775 & Lv8775));
assign Mzt775 = (~(Gwh675 | Eji675));
assign Yyt775 = (Tzt775 | Ye0775);
assign Bxt775 = (A0u775 & H0u775);
assign A0u775 = (~(O0u775 & Nxs775));
assign O0u775 = (~(Joi675 | Xhi675));
assign Nwt775 = (~(V0u775 | C1u775));
assign C1u775 = (Rpi675 ? J1u775 : Qf9775);
assign J1u775 = (Q1u775 & Aus775);
assign Q1u775 = (X1u775 & E2u775);
assign X1u775 = (~(L2u775 & S2u775));
assign L2u775 = (Z2u775 & G3u775);
assign G3u775 = (~(N3u775 & U3u775));
assign N3u775 = (~(Iq1775 | Jxj775));
assign Z2u775 = (~(Xhi675 & B4u775));
assign B4u775 = (~(I4u775 & P4u775));
assign P4u775 = (~(W4u775 | Ilk775));
assign I4u775 = (D5u775 & K5u775);
assign K5u775 = (Ia3775 | Qgi675);
assign D5u775 = (Jfi675 | Eji675);
assign V0u775 = (~(R5u775 & Y5u775));
assign Y5u775 = (~(Uo9775 & F6u775));
assign R5u775 = (~(Lv8775 & Ib9775));
assign Evt775 = (M6u775 & T6u775);
assign T6u775 = (A7u775 | U50775);
assign M6u775 = (Kls775 ? O7u775 : H7u775);
assign O7u775 = (~(V7u775 & Eh1775));
assign V7u775 = (Sh1775 & O4p675);
assign H7u775 = (~(C8u775 & A3k775));
assign C8u775 = (~(Ryf775 | Del775));
assign B0s675 = (!J8u775);
assign J8u775 = (hready_i ? Q8u775 : Zry675);
assign Q8u775 = (X8u775 & E9u775);
assign E9u775 = (L9u775 & S9u775);
assign S9u775 = (Z9u775 & Gau775);
assign Gau775 = (~(Nau775 & Uau775));
assign Uau775 = (Bbu775 | Ibu775);
assign Ibu775 = (Wk0775 & U50775);
assign Nau775 = (~(Vxo675 | Rto675));
assign Z9u775 = (~(Pbu775 | Lzb775));
assign Lzb775 = (My9775 & Ezo675);
assign Pbu775 = (Wbu775 & Qos775);
assign Wbu775 = (Jh0775 & Zck775);
assign L9u775 = (Dcu775 & Kcu775);
assign Kcu775 = (~(Rcu775 & Vsg775));
assign Rcu775 = (~(Nvg775 | Ycu775));
assign Dcu775 = (~(Srj775 & Fdu775));
assign Fdu775 = (~(Pw9775 & Mdu775));
assign Mdu775 = (Tdu775 | W1p675);
assign X8u775 = (Aeu775 & Heu775);
assign Heu775 = (Oeu775 & Veu775);
assign Veu775 = (Qsa775 | X7a775);
assign Oeu775 = (Cfu775 & Jfu775);
assign Jfu775 = (~(Qfu775 & Xza775));
assign Qfu775 = (~(Qsa775 & Xfu775));
assign Xfu775 = (~(My9775 & Egu775));
assign Egu775 = (~(Lgu775 & Sgu775));
assign Sgu775 = (~(Zgu775 & Zfa775));
assign Lgu775 = (~(Ghu775 & U50775));
assign Ghu775 = (Pw9775 | V8p675);
assign Qsa775 = (!Q7a775);
assign Q7a775 = (Lx6775 & X5p675);
assign Cfu775 = (~(Bbu775 & A3z675));
assign A3z675 = (~(Xuf775 | Xza775));
assign Aeu775 = (Nhu775 & Uhu775);
assign Uhu775 = (Biu775 | Vya775);
assign Nhu775 = (~(Iiu775 & E5z675));
assign Iiu775 = (~(Piu775 & Wiu775));
assign Wiu775 = (Dju775 & Kju775);
assign Kju775 = (Rju775 & Tst775);
assign Tst775 = (~(Yju775 & Fku775));
assign Yju775 = (~(Tsf775 | Wnb775));
assign Rju775 = (~(Mku775 | Rj9775));
assign Dju775 = (Tku775 & Alu775);
assign Alu775 = (~(Hlu775 & Vvr775));
assign Hlu775 = (Mwo675 & Olu775);
assign Olu775 = (K1z675 | T2r775);
assign Tku775 = (Vlu775 & Cmu775);
assign Vlu775 = (~(Jmu775 & Qmu775));
assign Qmu775 = (Frg775 & Ub1775);
assign Jmu775 = (~(Rba775 | I6l775));
assign Piu775 = (Xmu775 & Enu775);
assign Enu775 = (Lnu775 & Snu775);
assign Snu775 = (~(Eck775 & Zx6775));
assign Lnu775 = (Znu775 & Gou775);
assign Gou775 = (~(Nou775 & Uou775));
assign Nou775 = (~(M53775 | Lki675));
assign Znu775 = (~(Ous775 & Aus775));
assign Xmu775 = (~(Bpu775 | Ipu775));
assign Ipu775 = (Tli675 ? Ppu775 : Sta775);
assign Ppu775 = (~(A9l775 | Ahk775));
assign Bpu775 = (~(Wpu775 & Dqu775));
assign Dqu775 = (~(Rvb775 & T5a775));
assign Wpu775 = (Bvh675 ? Rqu775 : Kqu775);
assign Rqu775 = (Yqu775 & Fru775);
assign Fru775 = (Mru775 & Tru775);
assign Tru775 = (~(Gwh675 | V8p675));
assign Mru775 = (Asu775 & Hsu775);
assign Hsu775 = (~(Osu775 & Eji675));
assign Osu775 = (Qgi675 ? Ctu775 : Vsu775);
assign Ctu775 = (~(Jtu775 & Qtu775));
assign Qtu775 = (Ryt775 | On0775);
assign Jtu775 = (Tc3775 | Ye0775);
assign Vsu775 = (~(Ef3775 | Jfi675));
assign Asu775 = (~(Ous775 & Xtu775));
assign Xtu775 = (~(Euu775 & Tgk775));
assign Tgk775 = (~(Cei675 ^ Jfi675));
assign Euu775 = (~(Luu775 | X73775));
assign Yqu775 = (Suu775 & Zuu775);
assign Zuu775 = (Gvu775 | Ef3775);
assign Suu775 = (Nvu775 & Uvu775);
assign Uvu775 = (~(Bwu775 & Nc0775));
assign Bwu775 = (~(Iwu775 & Pwu775));
assign Pwu775 = (Ye0775 ? Nh9775 : Ef3775);
assign Iwu775 = (Wwu775 & Dxu775);
assign Dxu775 = (~(S2u775 & Luu775));
assign Wwu775 = (Eqk775 | Hk3775);
assign Nvu775 = (~(S2u775 & Hk3775));
assign Kqu775 = (Kxu775 & Rxu775);
assign Rxu775 = (~(Yxu775 & Kls775));
assign Yxu775 = (~(K7s775 | Ycu775));
assign Kxu775 = (Fyu775 | Nvg775);
assign Uzr675 = (Bct775 ? Iw1l85[0] : Myu775);
assign Myu775 = (~(Tyu775 & Azu775));
assign Azu775 = (Hzu775 & Ozu775);
assign Ozu775 = (~(Vzu775 & Xhi675));
assign Hzu775 = (~(C0v775 & Obi675));
assign Tyu775 = (Ict775 & J0v775);
assign J0v775 = (~(T7i675 & Q0v775));
assign Nzr675 = (~(X0v775 & E1v775));
assign E1v775 = (L1v775 & S1v775);
assign S1v775 = (~(Aft775 & Sy1l85[1]));
assign L1v775 = (Z1v775 & Oft775);
assign Z1v775 = (Vft775 | O02775);
assign O02775 = (G2v775 & N2v775);
assign N2v775 = (U2v775 & B3v775);
assign B3v775 = (~(I3v775 & P3v775));
assign U2v775 = (W3v775 & Ufb775);
assign W3v775 = (~(D4v775 & K4v775));
assign G2v775 = (R4v775 & Y4v775);
assign Y4v775 = (~(F5v775 & M5v775));
assign R4v775 = (Yhb775 | T5v775);
assign X0v775 = (A6v775 & H6v775);
assign H6v775 = (~(E52l85[0] & Ykt775));
assign A6v775 = (Fj3775 | O6v775);
assign Gzr675 = (!V6v775);
assign V6v775 = (hready_i ? C7v775 : Xza775);
assign C7v775 = (J7v775 & Q7v775);
assign Q7v775 = (X7v775 & E8v775);
assign E8v775 = (L8v775 & S8v775);
assign S8v775 = (~(Sry675 | Z8v775));
assign L8v775 = (Ky8775 & Sot775);
assign X7v775 = (G9v775 & N9v775);
assign N9v775 = (~(O4p675 & U9v775));
assign U9v775 = (~(Bav775 & Iav775));
assign Iav775 = (~(Pav775 & Srj775));
assign Pav775 = (~(Kls775 | Mwo675));
assign G9v775 = (Wav775 & Dbv775);
assign Dbv775 = (~(Tdg775 & Kbv775));
assign Kbv775 = (~(Rbv775 & Ybv775));
assign Ybv775 = (~(Fcv775 & Frg775));
assign Fcv775 = (~(Ycu775 | U50775));
assign Rbv775 = (~(Z8a775 & T5a775));
assign Wav775 = (~(Mcv775 & E2u775));
assign Mcv775 = (~(Tcv775 & Adv775));
assign Adv775 = (~(Hdv775 & Ik0775));
assign Hdv775 = (~(Oya775 | Ezo675));
assign Tcv775 = (~(Bbu775 & F3p675));
assign J7v775 = (Odv775 & Vdv775);
assign Vdv775 = (Cev775 & Jev775);
assign Jev775 = (Qev775 & Xev775);
assign Xev775 = (~(Bbu775 & Rcg775));
assign Bbu775 = (~(Q6b775 | Vya775));
assign Qev775 = (~(Efv775 & Vsg775));
assign Cev775 = (Lfv775 & Sfv775);
assign Sfv775 = (~(Zfv775 & Ggv775));
assign Ggv775 = (~(Ngv775 & Ugv775));
assign Ugv775 = (Bhv775 & Qt9775);
assign Bhv775 = (~(Bk0775 | Sta775));
assign Ngv775 = (Ihv775 & Phv775);
assign Phv775 = (Whv775 | Ye0775);
assign Ihv775 = (Div775 & Kiv775);
assign Kiv775 = (~(Riv775 & Jf9775));
assign Riv775 = (~(Xza775 | Zqi675));
assign Div775 = (~(Vtt775 & Obi675));
assign Lfv775 = (~(Yiv775 & E5z675));
assign Yiv775 = (~(Fjv775 & Mjv775));
assign Mjv775 = (Tjv775 & Akv775);
assign Akv775 = (Hkv775 & Okv775);
assign Okv775 = (~(Vkv775 & Efv775));
assign Vkv775 = (~(Clv775 | Fkg775));
assign Hkv775 = (~(Yqg775 | Jlv775));
assign Tjv775 = (Qlv775 & Xlv775);
assign Xlv775 = (~(Vvr775 & Emv775));
assign Emv775 = (~(Wdl775 & Lmv775));
assign Lmv775 = (~(Nzy675 & V0g775));
assign Qlv775 = (Smv775 & Zmv775);
assign Zmv775 = (~(Gnv775 & Mdg775));
assign Gnv775 = (~(Y1z675 | Bvh675));
assign Smv775 = (~(Nnv775 & Unv775));
assign Nnv775 = (~(U50775 | Jqh675));
assign Fjv775 = (Bov775 & Iov775);
assign Iov775 = (Pov775 & Wov775);
assign Wov775 = (~(Dpv775 & E2u775));
assign Dpv775 = (~(Kpv775 & Rpv775));
assign Rpv775 = (Ypv775 & Fqv775);
assign Fqv775 = (~(Bk0775 & Mqv775));
assign Mqv775 = (~(Tqv775 & Arv775));
assign Arv775 = (Hrv775 & Orv775);
assign Hrv775 = (~(Xhi675 & Vrv775));
assign Vrv775 = (Nh9775 | Ilk775);
assign Tqv775 = (Csv775 & Jsv775);
assign Jsv775 = (Iq1775 | Eji675);
assign Csv775 = (Ia3775 ? Lyj775 : Ogs775);
assign Ypv775 = (~(Mku775 | Qsv775));
assign Mku775 = (Dia775 & Nc0775);
assign Dia775 = (Aus775 & Tli675);
assign Kpv775 = (Xsv775 & Etv775);
assign Etv775 = (~(Dqg775 & Sta775));
assign Xsv775 = (~(W4u775 & Gw8775));
assign Pov775 = (Ltv775 & Stv775);
assign Stv775 = (~(Z8a775 & Ztv775));
assign Ztv775 = (~(O4p675 & Guv775));
assign Guv775 = (R1z675 | Kls775);
assign Ltv775 = (~(Jf9775 & Nuv775));
assign Nuv775 = (~(Uuv775 & Bvv775));
assign Bvv775 = (Ryt775 | Ezo675);
assign Uuv775 = (Ivv775 & U50775);
assign Ivv775 = (~(Pvv775 & J7p675));
assign Pvv775 = (~(P58775 | F3p675));
assign Bov775 = (Wvv775 & Dwv775);
assign Dwv775 = (~(Nxs775 & Kwv775));
assign Kwv775 = (~(Rwv775 & Ywv775));
assign Ywv775 = (~(Bni675 & Fxv775));
assign Fxv775 = (~(Mxv775 & Txv775));
assign Txv775 = (~(Izk775 ^ Xhi675));
assign Mxv775 = (Ayv775 & Hyv775);
assign Hyv775 = (A9l775 | Tc3775);
assign Ayv775 = (Lyj775 | Lki675);
assign Rwv775 = (Oyv775 & Vyv775);
assign Vyv775 = (~(Czv775 & Joi675));
assign Czv775 = (Xhi675 & Jzv775);
assign Jzv775 = (~(Yzs775 & Qzv775));
assign Qzv775 = (~(Xzv775 & Iw2775));
assign Oyv775 = (~(E0w775 & Tc3775));
assign E0w775 = (~(L0w775 & Ia3775));
assign L0w775 = (~(Qgi675 ^ Eji675));
assign Wvv775 = (~(Rj9775 & M53775));
assign Odv775 = (S0w775 & O5b775);
assign S0w775 = (Z0w775 & G1w775);
assign G1w775 = (M7t775 | Dj9775);
assign Z0w775 = (Za1775 | Zfh775);
assign Zyr675 = (!N1w775);
assign N1w775 = (hready_i ? U1w775 : U50775);
assign U1w775 = (B2w775 & I2w775);
assign I2w775 = (P2w775 & W2w775);
assign W2w775 = (D3w775 & K3w775);
assign K3w775 = (R3w775 & Y3w775);
assign R3w775 = (Ugh775 & Sot775);
assign Sot775 = (Oya775 | F4w775);
assign Ugh775 = (~(Dba775 & M4w775));
assign D3w775 = (T4w775 & A5w775);
assign A5w775 = (~(H5w775 & Qnt775));
assign Qnt775 = (~(Oya775 | Ycu775));
assign H5w775 = (Ria775 & Ik0775);
assign T4w775 = (~(O5w775 & V5w775));
assign V5w775 = (~(Af1775 | Gwh675));
assign O5w775 = (S2u775 & Zfv775);
assign P2w775 = (C6w775 & J6w775);
assign J6w775 = (Q6w775 & X6w775);
assign X6w775 = (~(E7w775 & Vwj775));
assign E7w775 = (Xhi675 ? S7w775 : L7w775);
assign S7w775 = (~(Z7w775 & P5t775));
assign P5t775 = (!Pds775);
assign Pds775 = (Eji675 & Ilk775);
assign Z7w775 = (Gvu775 | Qgi675);
assign L7w775 = (Ogs775 & W4u775);
assign Q6w775 = (~(Yuj775 & G8w775));
assign G8w775 = (~(Cm9775 & N8w775));
assign N8w775 = (~(Tli675 & U8w775));
assign U8w775 = (~(Tzt775 & B9w775));
assign B9w775 = (~(Vjb775 & Eji675));
assign Cm9775 = (!Qsv775);
assign Qsv775 = (I9w775 & Tc3775);
assign C6w775 = (P9w775 & W9w775);
assign W9w775 = (~(Ub1775 & Daw775));
assign Daw775 = (~(M2k775 & Kaw775));
assign Kaw775 = (~(Raw775 & D3b775));
assign Raw775 = (~(I6l775 | Yaw775));
assign P9w775 = (~(Vsg775 & Fbw775));
assign Fbw775 = (~(Mbw775 & Tbw775));
assign Tbw775 = (Za1775 | Ycu775);
assign B2w775 = (Acw775 & Hcw775);
assign Hcw775 = (Ocw775 & Vcw775);
assign Vcw775 = (Cdw775 & Jdw775);
assign Jdw775 = (Bav775 | F3p675);
assign Cdw775 = (Qdw775 & Xdw775);
assign Xdw775 = (~(Eew775 & Lew775));
assign Lew775 = (~(Sew775 & Zew775));
assign Zew775 = (~(Gfw775 & T17775));
assign Gfw775 = (~(Nfw775 & Ufw775));
assign Ufw775 = (Bgw775 & Biu775);
assign Biu775 = (~(Igw775 & V8p675));
assign Igw775 = (~(D1z675 | Ezo675));
assign Bgw775 = (~(Pgw775 & Jf9775));
assign Pgw775 = (Wgw775 & Y1z675);
assign Wgw775 = (~(Dhw775 & Khw775));
assign Khw775 = (Hk3775 | Gwh675);
assign Nfw775 = (Rhw775 & Yhw775);
assign Yhw775 = (~(Pxf775 & V8p675));
assign Rhw775 = (Q6b775 | F3p675);
assign Sew775 = (~(Fiw775 & Xt2775));
assign Qdw775 = (~(S8a775 & Miw775));
assign Ocw775 = (Tiw775 & Ajw775);
assign Ajw775 = (~(Hjw775 & Lis775));
assign Lis775 = (~(Ep0775 & Ojw775));
assign Ojw775 = (~(Wk0775 & M7t775));
assign Tiw775 = (~(Vjw775 & E5z675));
assign Vjw775 = (~(Ckw775 & Jkw775));
assign Jkw775 = (Pub775 & Qkw775);
assign Pub775 = (~(Vtt775 & Xza775));
assign Ckw775 = (Xkw775 & Elw775);
assign Elw775 = (~(Rvb775 & Iah775));
assign Xkw775 = (~(Llw775 & Iek775));
assign Acw775 = (Slw775 & Zlw775);
assign Zlw775 = (Gmw775 & Nmw775);
assign Nmw775 = (~(Bni675 & Umw775));
assign Umw775 = (~(Bnw775 & Inw775));
assign Inw775 = (Pnw775 & Wnw775);
assign Wnw775 = (~(Dow775 & Kow775));
assign Kow775 = (Row775 & M71775);
assign Row775 = (~(Yow775 & Fpw775));
assign Fpw775 = (~(Mpw775 & Eji675));
assign Yow775 = (Eqk775 | M53775);
assign Dow775 = (Uo9775 & Zfv775);
assign Pnw775 = (Tpw775 | Chs775);
assign Chs775 = (~(Xzv775 & Cei675));
assign Xzv775 = (~(Jfi675 | Qgi675));
assign Tpw775 = (~(Vgs775 & Vci675));
assign Bnw775 = (Aqw775 & Hqw775);
assign Hqw775 = (~(Xxj775 & Oqw775));
assign Oqw775 = (~(Qgi675 & Vqw775));
assign Vqw775 = (Tc3775 | On0775);
assign Aqw775 = (~(Yuj775 & C89775));
assign Gmw775 = (~(Vvr775 & Crw775));
assign Crw775 = (~(Jrw775 & Qrw775));
assign Qrw775 = (Xrw775 & Esw775);
assign Esw775 = (~(Lsw775 & Ssw775));
assign Ssw775 = (~(K7s775 & Fyu775));
assign Xrw775 = (Zsw775 & Gtw775);
assign Gtw775 = (~(Ntw775 & Utw775));
assign Ntw775 = (~(Dwa775 | Wxf775));
assign Zsw775 = (~(Buw775 & F6g775));
assign Buw775 = (~(Q91775 | Lrh675));
assign Jrw775 = (Iuw775 & Puw775);
assign Puw775 = (~(Lh1775 & Wuw775));
assign Wuw775 = (~(U3g775 & Dvw775));
assign Dvw775 = (~(Kvw775 & Xza775));
assign Kvw775 = (Pw9775 | P58775);
assign Iuw775 = (~(Rvw775 & T17775));
assign Rvw775 = (~(Yvw775 & Fww775));
assign Fww775 = (~(Mww775 & Zfv775));
assign Mww775 = (~(Pw9775 | Rto675));
assign Yvw775 = (F4w775 | Xuf775);
assign Slw775 = (~(Tww775 | Axw775));
assign Axw775 = (~(Te1775 | Fkg775));
assign Tww775 = (O4p675 ? Hxw775 : Qza775);
assign Hxw775 = (~(Oxw775 & Vxw775));
assign Vxw775 = (L2g775 | Eta775);
assign Oxw775 = (Cyw775 & Jyw775);
assign Jyw775 = (~(Miw775 & Fvq775));
assign Cyw775 = (~(Lps775 & Rba775));
assign Syr675 = (~(Qyw775 & Xyw775));
assign Xyw775 = (~(X5p675 & Ezw775));
assign Ezw775 = (~(Lzw775 & hready_i));
assign Lzw775 = (~(Szw775 | Hjw775));
assign Szw775 = (~(V8p675 | W1p675));
assign Qyw775 = (~(hready_i & Zzw775));
assign Zzw775 = (~(G0x775 & N0x775));
assign N0x775 = (U0x775 & B1x775);
assign B1x775 = (~(Wnb775 & I1x775));
assign I1x775 = (~(P1x775 & W1x775));
assign W1x775 = (~(D2x775 & Z8a775));
assign D2x775 = (~(Vxo675 | O4p675));
assign P1x775 = (Tsf775 | Wxf775);
assign Tsf775 = (!Rvb775);
assign U0x775 = (K2x775 & Dj9775);
assign K2x775 = (~(R2x775 & Gwh675));
assign R2x775 = (Rpi675 & Y2x775);
assign Y2x775 = (~(Af1775 & F3x775));
assign F3x775 = (~(M3x775 & O0g775));
assign O0g775 = (N0p675 & Cg8775);
assign G0x775 = (T3x775 & A4x775);
assign A4x775 = (Te1775 | E5z675);
assign T3x775 = (O3k775 & H4x775);
assign H4x775 = (B0z675 | Xxq775);
assign O3k775 = (~(Dba775 & Zx6775));
assign Lyr675 = (A27775 ? Ceh775 : J7p675);
assign Eyr675 = (~(O4x775 & V4x775));
assign V4x775 = (C5x775 | J5x775);
assign O4x775 = (X5x775 ? N1p775 : Q5x775);
assign Q5x775 = (E6x775 & L6x775);
assign L6x775 = (S6x775 & Z6x775);
assign Z6x775 = (Pi9775 & Dj9775);
assign Pi9775 = (~(Per775 & X5p675));
assign S6x775 = (G7x775 & N7x775);
assign N7x775 = (~(U7x775 & Lki675));
assign U7x775 = (B8x775 & Nc0775);
assign B8x775 = (~(Wva775 & I8x775));
assign I8x775 = (~(N9a775 & Zfv775));
assign Wva775 = (Lws775 | Lrh675);
assign Lws775 = (!I9w775);
assign I9w775 = (Ous775 & Bvh675);
assign G7x775 = (~(P8x775 & Nfn675));
assign E6x775 = (W8x775 & D9x775);
assign D9x775 = (Xt2775 | K9x775);
assign W8x775 = (R9x775 & Y9x775);
assign Y9x775 = (Iw2775 | Fax775);
assign R9x775 = (~(Kr1775 & Eji675));
assign Xxr675 = (!Max775);
assign Max775 = (hready_i ? Tax775 : Wks775);
assign Tax775 = (Abx775 & Hbx775);
assign Hbx775 = (~(Obx775 & Vbx775));
assign Qxr675 = (!Ccx775);
assign Ccx775 = (hready_i ? Jcx775 : Y1z675);
assign Jcx775 = (Qcx775 & Xcx775);
assign Xcx775 = (Edx775 & Ldx775);
assign Ldx775 = (Sdx775 & Zdx775);
assign Zdx775 = (Qkw775 & Jrb775);
assign Qkw775 = (~(Gex775 & Fiw775));
assign Gex775 = (~(Q91775 | Rto675));
assign Sdx775 = (Ggh775 & Nex775);
assign Edx775 = (Uex775 & Bfx775);
assign Bfx775 = (~(Ifx775 & Iso675));
assign Ifx775 = (~(B0z675 | Za1775));
assign Uex775 = (Pfx775 & Y3w775);
assign Pfx775 = (~(Wfx775 & Iek775));
assign Wfx775 = (~(Pb9775 | Kq9775));
assign Kq9775 = (Tli675 & Rpi675);
assign Qcx775 = (Dgx775 & Kgx775);
assign Kgx775 = (Rgx775 & Ygx775);
assign Ygx775 = (~(Eh1775 & D7l775));
assign Rgx775 = (Fhx775 & Mhx775);
assign Mhx775 = (~(Thx775 & Zry675));
assign Thx775 = (~(Aix775 & Hix775));
assign Hix775 = (Veg775 | Cg8775);
assign Aix775 = (Oix775 & Vix775);
assign Vix775 = (~(Zgu775 & Zsb775));
assign Zgu775 = (~(E5z675 | Kls775));
assign Oix775 = (Wks775 | B2b775);
assign Fhx775 = (~(Cjx775 & M71775));
assign Cjx775 = (~(Jjx775 & Qjx775));
assign Qjx775 = (Xjx775 & Ekx775);
assign Ekx775 = (Lkx775 & Skx775);
assign Skx775 = (~(Zkx775 & Mvj775));
assign Zkx775 = (Glx775 & E2u775);
assign Glx775 = (~(Nlx775 & Ulx775));
assign Ulx775 = (~(Bmx775 & Tc3775));
assign Bmx775 = (~(Imx775 & U4t775));
assign U4t775 = (Pmx775 & Wmx775);
assign Wmx775 = (~(Dnx775 & Eji675));
assign Dnx775 = (~(Iq1775 | Xhi675));
assign Pmx775 = (~(Lki675 & Knx775));
assign Knx775 = (Xhi675 | Ogs775);
assign Imx775 = (Rpi675 & Rnx775);
assign Rnx775 = (A9l775 | Lyj775);
assign Nlx775 = (~(Kzs775 & Dqg775));
assign Lkx775 = (~(Ynx775 & Tli675));
assign Ynx775 = (Joi675 & Fox775);
assign Fox775 = (~(Mox775 & Tox775));
assign Tox775 = (~(Apx775 & Hpx775));
assign Hpx775 = (Opx775 & Jxj775);
assign Jxj775 = (Xhi675 & On0775);
assign Opx775 = (Izk775 & Nxs775);
assign Apx775 = (Vpx775 & Cqx775);
assign Vpx775 = (Jpk775 & Yzs775);
assign Mox775 = (Tzt775 | Jqx775);
assign Xjx775 = (Qqx775 & Xqx775);
assign Xqx775 = (~(Erx775 & Cqx775));
assign Erx775 = (W4u775 & Uo9775);
assign Qqx775 = (~(Efv775 & Rvb775));
assign Efv775 = (~(Te1775 | Kls775));
assign Jjx775 = (Lrx775 & Srx775);
assign Srx775 = (Zrx775 & Gsx775);
assign Gsx775 = (~(Nsx775 & Cut775));
assign Zrx775 = (~(Ib9775 & Usx775));
assign Usx775 = (~(Btx775 & Itx775));
assign Btx775 = (Ptx775 & Wtx775);
assign Wtx775 = (~(Dux775 & Sta775));
assign Dux775 = (Tc3775 ? X73775 : U3u775);
assign Ptx775 = (~(Gw8775 & Izk775));
assign Lrx775 = (Of1775 & Kux775);
assign Kux775 = (~(S2u775 & Uou775));
assign Of1775 = (Rux775 | Za1775);
assign Dgx775 = (Yux775 & Fvx775);
assign Fvx775 = (W1p675 ? Tvx775 : Mvx775);
assign Tvx775 = (~(N0p675 & Awx775));
assign Awx775 = (~(Fkg775 & Ndk775));
assign Ndk775 = (E5z675 | Eta775);
assign Mvx775 = (~(Dba775 & Xza775));
assign Yux775 = (Ct9775 & Hwx775);
assign Hwx775 = (Kba775 | O4p675);
assign Kba775 = (!Osg775);
assign Jxr675 = (Owx775 & Vwx775);
assign Vwx775 = (~(Cxx775 & Jxx775));
assign Jxx775 = (Qxx775 & Xxx775);
assign Xxx775 = (Eyx775 & Lyx775);
assign Lyx775 = (Syx775 & Zyx775);
assign Syx775 = (~(Gzx775 & Vgs775));
assign Vgs775 = (Nzx775 & Uzx775);
assign Uzx775 = (~(B0y775 | M53775));
assign B0y775 = (!Dc9775);
assign Dc9775 = (Izk775 & Tli675);
assign Nzx775 = (Yzs775 & Ncs775);
assign Ncs775 = (!I0y775);
assign Yzs775 = (P0y775 & Ora775);
assign P0y775 = (~(Hai675 | Obi675));
assign Gzx775 = (Jpk775 & W0y775);
assign W0y775 = (Iw2775 | On0775);
assign Jpk775 = (~(Cei675 | Qgi675));
assign Eyx775 = (D1y775 & K1y775);
assign K1y775 = (~(R1y775 & Uo9775));
assign R1y775 = (Wc1775 & Y1y775);
assign Y1y775 = (~(F2y775 & M2y775));
assign M2y775 = (~(T2y775 & Mpw775));
assign T2y775 = (~(X73775 | Ye0775));
assign F2y775 = (Hk3775 | Ef3775);
assign D1y775 = (~(A3y775 & Iek775));
assign A3y775 = (H3y775 & E5z675);
assign H3y775 = (~(Itx775 & O3y775));
assign O3y775 = (~(V3y775 & Dqg775));
assign Dqg775 = (Ia3775 & Tc3775);
assign V3y775 = (~(Ahk775 | Xhi675));
assign Itx775 = (C4y775 | Ye0775);
assign Qxx775 = (J4y775 & Q4y775);
assign Q4y775 = (X4y775 & E5y775);
assign E5y775 = (~(L5y775 & M3x775));
assign L5y775 = (~(Eot775 | Oya775));
assign X4y775 = (~(S5y775 & Z5y775));
assign S5y775 = (~(Za1775 | N0p675));
assign J4y775 = (G6y775 & N6y775);
assign N6y775 = (~(U6y775 & Gjs775));
assign U6y775 = (~(K7s775 | Y1z675));
assign G6y775 = (~(Xxq775 & B7y775));
assign B7y775 = (Osg775 | Gjs775);
assign Cxx775 = (I7y775 & P7y775);
assign P7y775 = (W7y775 & D8y775);
assign D8y775 = (K8y775 & R8y775);
assign R8y775 = (~(T5a775 & Y8y775));
assign Y8y775 = (~(F9y775 & M9y775));
assign M9y775 = (~(Dba775 & N0p675));
assign F9y775 = (~(A3k775 & W1p675));
assign K8y775 = (~(Bsk775 & Zfv775));
assign Bsk775 = (Utw775 & Nsx775);
assign Utw775 = (T9y775 & Aay775);
assign T9y775 = (Hay775 & Oay775);
assign W7y775 = (Vay775 & Cby775);
assign Cby775 = (~(Kls775 & Jby775));
assign Jby775 = (~(Qby775 & Xby775));
assign Xby775 = (~(A3k775 & Ecy775));
assign Ecy775 = (S8a775 | Lcy775);
assign Lcy775 = (Zfa775 & Q91775);
assign S8a775 = (Zx6775 & W1p675);
assign Qby775 = (Scy775 & Zcy775);
assign Zcy775 = (~(Gdy775 & Ndy775));
assign Ndy775 = (~(Ep0775 | Rto675));
assign Gdy775 = (Qos775 & Mdg775);
assign Mdg775 = (Nzy675 & Zry675);
assign Scy775 = (~(Udy775 & C1g775));
assign Udy775 = (Frg775 & E5z675);
assign Vay775 = (~(Bey775 & M71775));
assign Bey775 = (~(Iey775 & Pey775));
assign Pey775 = (Wey775 & Sng775);
assign Sng775 = (~(Dfy775 & Ik0775));
assign Dfy775 = (Rj9775 & Gvu775);
assign Wey775 = (~(Kfy775 & Rfy775));
assign Rfy775 = (~(Tli675 | Rpi675));
assign Kfy775 = (U2a775 & E2u775);
assign Iey775 = (Yfy775 & Fgy775);
assign Fgy775 = (~(Mgy775 & Ik0775));
assign Mgy775 = (Rj9775 & Xhi675);
assign Yfy775 = (Fkg775 | Pw9775);
assign I7y775 = (Tgy775 & Ahy775);
assign Ahy775 = (~(Wsk775 | Q4k775));
assign Q4k775 = (~(Hhy775 & Ohy775));
assign Ohy775 = (~(Jh0775 & Xza775));
assign Jh0775 = (Rvb775 & Tdg775);
assign Hhy775 = (Crb775 & Vhy775);
assign Crb775 = (~(Hjw775 & Dba775));
assign Wsk775 = (~(Ciy775 & hready_i));
assign Ciy775 = (Y3w775 & Nb1775);
assign Nb1775 = (!Jiy775);
assign Tgy775 = (Qiy775 & Zps775);
assign Zps775 = (Xiy775 & Ejy775);
assign Ejy775 = (~(Xxj775 & Lyj775));
assign Xxj775 = (~(I0y775 | Orv775));
assign Xiy775 = (Ljy775 & Sjy775);
assign Sjy775 = (~(Zjy775 & Gjs775));
assign Gjs775 = (Tdg775 & Vvr775);
assign Zjy775 = (~(W1p675 | F3p675));
assign Ljy775 = (I0y775 | Bni675);
assign I0y775 = (~(Iek775 & Q89775));
assign Iek775 = (~(Nc0775 | V8p675));
assign Qiy775 = (Rpi675 ? Nky775 : Gky775);
assign Nky775 = (~(Vwj775 & Uky775));
assign Uky775 = (~(Bly775 & Ily775));
assign Ily775 = (Qgi675 ? Wly775 : Ply775);
assign Wly775 = (Kzs775 | Lki675);
assign Bly775 = (Dmy775 & A9l775);
assign A9l775 = (!Owj775);
assign Dmy775 = (~(Ogs775 & Xpk775));
assign Ogs775 = (Kmy775 & Rpa775);
assign Rpa775 = (T7i675 & A9i675);
assign Kmy775 = (~(Mr2775 | Iq1775));
assign Mr2775 = (!Hai675);
assign Vwj775 = (Rmy775 & Yuj775);
assign Rmy775 = (~(C4y775 | Joi675));
assign Gky775 = (~(Ymy775 & Yuj775));
assign Yuj775 = (~(Jqx775 | Yaw775));
assign Ymy775 = (Tli675 & Fny775);
assign Fny775 = (~(Pb9775 & Mny775));
assign Mny775 = (~(Owj775 & N9a775));
assign Owj775 = (Ia3775 & X73775);
assign Pb9775 = (!Mvj775);
assign Owx775 = (N0p675 | hready_i);
assign Cxr675 = (Tny775 & Aoy775);
assign Aoy775 = (~(Hoy775 & Ooy775));
assign Ooy775 = (Voy775 & Cpy775);
assign Cpy775 = (Jpy775 & Qpy775);
assign Qpy775 = (Xpy775 & Eqy775);
assign Eqy775 = (~(Ous775 & Lqy775));
assign Lqy775 = (~(C4y775 & Sqy775));
assign Sqy775 = (~(Nxs775 & Zqy775));
assign Zqy775 = (~(Gry775 & Nry775));
assign Nry775 = (Ury775 & Ia3775);
assign Ury775 = (Vci675 | Jfi675);
assign Gry775 = (~(Iq1775 | Ty2775));
assign Xpy775 = (~(C89775 & Bsy775));
assign Bsy775 = (~(Isy775 & Psy775));
assign Psy775 = (~(Cqx775 & Wsy775));
assign Wsy775 = (~(Dty775 & Kty775));
assign Kty775 = (Tc3775 | Jfi675);
assign Dty775 = (~(Ilk775 | Xhi675));
assign Isy775 = (~(Ria775 & Nh9775));
assign Jpy775 = (Rty775 & Yty775);
assign Yty775 = (~(Z8a775 & Fuy775));
assign Fuy775 = (~(Muy775 & Tuy775));
assign Tuy775 = (~(Avy775 & Hvy775));
assign Hvy775 = (Ovy775 & Rba775);
assign Ovy775 = (Sh1775 | Ex6775);
assign Ex6775 = (F3p675 & Zry675);
assign Muy775 = (~(Hjw775 & M7t775));
assign Hjw775 = (Zry675 & D1z675);
assign Rty775 = (~(Kls775 & Vvy775));
assign Vvy775 = (~(Cwy775 & Jwy775));
assign Jwy775 = (~(Qwy775 & Frg775));
assign Qwy775 = (~(U3g775 | F3p675));
assign Cwy775 = (~(Eck775 & Fvq775));
assign Voy775 = (Xwy775 & Exy775);
assign Exy775 = (Lxy775 & Sxy775);
assign Sxy775 = (~(Zxy775 & Cm2775));
assign Zxy775 = (~(Gyy775 & Nyy775));
assign Nyy775 = (Agl775 | O4p675);
assign Gyy775 = (~(C1g775 & Nzy675));
assign Lxy775 = (~(Vtt775 & Cg8775));
assign Xwy775 = (Uyy775 & Bzy775);
assign Bzy775 = (Att775 | Lrh675);
assign Uyy775 = (~(Vvr775 & Izy775));
assign Izy775 = (~(Pzy775 & Wzy775));
assign Wzy775 = (L2g775 | Q91775);
assign Pzy775 = (D0z775 & K0z775);
assign K0z775 = (I6l775 | Rto675);
assign D0z775 = (A2l775 | Xuf775);
assign Hoy775 = (R0z775 & Y0z775);
assign Y0z775 = (F1z775 & M1z775);
assign M1z775 = (T1z775 & A2z775);
assign A2z775 = (~(Rpi675 & H2z775));
assign H2z775 = (~(O2z775 & V2z775));
assign V2z775 = (Eqk775 | J6b775);
assign O2z775 = (C3z775 & J3z775);
assign J3z775 = (~(Q3z775 & Ria775));
assign Q3z775 = (~(Cm2775 | Xhi675));
assign C3z775 = (~(D6t775 & Nxs775));
assign T1z775 = (~(Rvb775 & X3z775));
assign X3z775 = (E4z775 | L4z775);
assign L4z775 = (Mwo675 ? K1z675 : Kny675);
assign E4z775 = (~(S4z775 & Fyu775));
assign Fyu775 = (Wnb775 | Vxo675);
assign S4z775 = (Te1775 | Qos775);
assign F1z775 = (Z4z775 & G5z775);
assign G5z775 = (~(N5z775 & Nc0775));
assign N5z775 = (~(U5z775 & B6z775));
assign B6z775 = (I6z775 & P6z775);
assign P6z775 = (~(Gw8775 & Lki675));
assign I6z775 = (W6z775 & D7z775);
assign D7z775 = (~(K7z775 & Cqx775));
assign K7z775 = (~(Cm2775 | U3u775));
assign W6z775 = (~(Bk0775 & R7z775));
assign R7z775 = (~(Y7z775 & F8z775));
assign F8z775 = (X73775 ? Wp9775 : Jfi675);
assign Wp9775 = (!Ilk775);
assign Y7z775 = (~(Kzs775 | Fgk775));
assign Kzs775 = (On0775 & M53775);
assign U5z775 = (M8z775 & T8z775);
assign T8z775 = (~(Vjb775 & Tc3775));
assign Vjb775 = (Bvh675 & Hk3775);
assign M8z775 = (Ahk775 | Rpi675);
assign Z4z775 = (~(Jf9775 & Psk775));
assign R0z775 = (~(A9z775 | H9z775));
assign H9z775 = (W1p675 ? O9z775 : Jiy775);
assign O9z775 = (Fyg775 & Bek775);
assign Bek775 = (~(Wks775 & E5z675));
assign Jiy775 = (Unv775 & N0p675);
assign A9z775 = (V9z775 | H8t775);
assign H8t775 = (~(Caz775 & Jaz775));
assign Jaz775 = (Qaz775 & Xaz775);
assign Xaz775 = (~(Ebz775 & V8p675));
assign Ebz775 = (~(Pw9775 | W1p675));
assign Qaz775 = (Qt9775 & Jrb775);
assign Qt9775 = (!Qf9775);
assign Qf9775 = (Gwh675 & Bvh675);
assign Caz775 = (hready_i & Lbz775);
assign V9z775 = (Tli675 ? Sbz775 : Rj9775);
assign Tny775 = (Mwo675 | hready_i);
assign Vwr675 = (Zbz775 | Gcz775);
assign Gcz775 = (~(Ncz775 | J5x775));
assign Zbz775 = (X5x775 ? Byi675 : Ucz775);
assign Ucz775 = (~(Bdz775 & Idz775));
assign Idz775 = (Pdz775 & Wdz775);
assign Wdz775 = (~(P8x775 & Xgn675));
assign P8x775 = (P8n675 & Dez775);
assign Dez775 = (~(Kez775 & Lvf775));
assign Kez775 = (~(Ddt775 | Qza775));
assign Pdz775 = (Ty2775 | Fax775);
assign Bdz775 = (Rez775 & Yez775);
assign Yez775 = (~(Kr1775 & Lki675));
assign Kr1775 = (Sbz775 & Zfv775);
assign Rez775 = (Iw2775 | K9x775);
assign Owr675 = (!Ffz775);
assign Ffz775 = (A27775 ? M2s675 : X7a775);
assign A27775 = (~(Lcz675 | Cg8775));
assign M2s675 = (~(P8n675 & Mfz775));
assign Mfz775 = (~(Tfz775 & Agz775));
assign Agz775 = (Hgz775 & Ogz775);
assign Ogz775 = (~(Bln675 | Lmn675));
assign Hgz775 = (~(Hin675 | Rjn675));
assign Tfz775 = (Vgz775 & Chz775);
assign Chz775 = (~(Rqn675 | Csn675));
assign Vgz775 = (~(Vnn675 | Gpn675));
assign Hwr675 = (~(Jhz775 & Qhz775));
assign Qhz775 = (Xhz775 & Eiz775);
assign Eiz775 = (~(E52l85[21] & Ykt775));
assign Xhz775 = (Liz775 & Siz775);
assign Siz775 = (Vft775 | D8d775);
assign D8d775 = (Ziz775 & Gjz775);
assign Gjz775 = (Njz775 & Ujz775);
assign Ujz775 = (~(Bkz775 & Dkt775));
assign Njz775 = (Ikz775 | Nit775);
assign Ziz775 = (Pkz775 & Wkz775);
assign Wkz775 = (~(Pjt775 & Dlz775));
assign Pkz775 = (~(Lht775 & Klz775));
assign Liz775 = (~(Aft775 & Sy1l85[22]));
assign Jhz775 = (Rlz775 & Ylz775);
assign Ylz775 = (~(vis_pc_o[21] & P60775));
assign Awr675 = (~(Fmz775 & Mmz775));
assign Mmz775 = (Tmz775 & Anz775);
assign Anz775 = (~(Aft775 & Sy1l85[31]));
assign Tmz775 = (Hnz775 & Oft775);
assign Hnz775 = (Vft775 | B1c775);
assign B1c775 = (Onz775 & Vnz775);
assign Vnz775 = (Coz775 & Joz775);
assign Joz775 = (~(Qoz775 & Wjt775));
assign Coz775 = (Xoz775 & Zht775);
assign Xoz775 = (Git775 | Epz775);
assign Onz775 = (Lpz775 & Spz775);
assign Spz775 = (~(Zpz775 & Eht775));
assign Lpz775 = (Gqz775 | Nqz775);
assign Fmz775 = (Uqz775 & Brz775);
assign Brz775 = (~(E52l85[30] & Ykt775));
assign Uqz775 = (~(vis_pc_o[30] & P60775));
assign Tvr675 = (Lcz675 ? Plo675 : Irz775);
assign Irz775 = (!Prz775);
assign Mvr675 = (Jm2775 ? Eko675 : Ndz675);
assign Fvr675 = (~(Wrz775 & Dsz775));
assign Dsz775 = (~(Ksz775 & hrdata_i[16]));
assign Wrz775 = (~(Uxn675 & Jm2775));
assign Yur675 = (~(Rsz775 & Ysz775));
assign Ysz775 = (~(Ksz775 & hrdata_i[17]));
assign Rsz775 = (~(Ezn675 & Jm2775));
assign Rur675 = (~(Ftz775 & Mtz775));
assign Mtz775 = (~(Ksz775 & hrdata_i[18]));
assign Ftz775 = (~(O0o675 & Jm2775));
assign Kur675 = (~(Ttz775 & Auz775));
assign Auz775 = (~(Ksz775 & hrdata_i[19]));
assign Ttz775 = (~(Y1o675 & Jm2775));
assign Dur675 = (~(Huz775 & Ouz775));
assign Ouz775 = (~(Ksz775 & hrdata_i[20]));
assign Huz775 = (~(I3o675 & Jm2775));
assign Wtr675 = (~(Vuz775 & Cvz775));
assign Cvz775 = (~(Ksz775 & hrdata_i[21]));
assign Vuz775 = (~(S4o675 & Jm2775));
assign Ptr675 = (~(Jvz775 & Qvz775));
assign Qvz775 = (~(Ksz775 & hrdata_i[22]));
assign Jvz775 = (~(C6o675 & Jm2775));
assign Itr675 = (~(Xvz775 & Ewz775));
assign Ewz775 = (~(Ksz775 & hrdata_i[23]));
assign Xvz775 = (~(M7o675 & Jm2775));
assign Btr675 = (~(Lwz775 & Swz775));
assign Swz775 = (~(Ksz775 & hrdata_i[24]));
assign Lwz775 = (~(W8o675 & Jm2775));
assign Usr675 = (~(Zwz775 & Gxz775));
assign Gxz775 = (~(Ksz775 & hrdata_i[25]));
assign Zwz775 = (~(Gao675 & Jm2775));
assign Nsr675 = (~(Nxz775 & Uxz775));
assign Uxz775 = (~(Ksz775 & hrdata_i[26]));
assign Nxz775 = (~(Qbo675 & Jm2775));
assign Gsr675 = (~(Byz775 & Iyz775));
assign Iyz775 = (~(Ksz775 & hrdata_i[27]));
assign Byz775 = (~(Bdo675 & Jm2775));
assign Zrr675 = (~(Pyz775 & Wyz775));
assign Wyz775 = (~(Ksz775 & hrdata_i[28]));
assign Pyz775 = (~(Meo675 & Jm2775));
assign Srr675 = (~(Dzz775 & Kzz775));
assign Kzz775 = (~(Ksz775 & hrdata_i[29]));
assign Dzz775 = (~(Xfo675 & Jm2775));
assign Lrr675 = (~(Rzz775 & Yzz775));
assign Yzz775 = (~(Ksz775 & hrdata_i[30]));
assign Rzz775 = (~(Iho675 & Jm2775));
assign Err675 = (~(F00875 & M00875));
assign M00875 = (~(Ksz775 & hrdata_i[31]));
assign Ksz775 = (~(Ndz675 | Jm2775));
assign Ndz675 = (!Kfz675);
assign Kfz675 = (T00875 & vis_tbit_o);
assign T00875 = (~(hresp_i | Zmo675));
assign F00875 = (~(Tio675 & Jm2775));
assign Jm2775 = (!Nn3775);
assign Nn3775 = (Plo675 & hready_i);
assign Xqr675 = (Bct775 ? Iw1l85[1] : A10875);
assign A10875 = (~(H10875 & O10875));
assign O10875 = (V10875 & C20875);
assign C20875 = (~(C0v775 & Vci675));
assign V10875 = (J20875 & Q20875);
assign Q20875 = (~(X20875 & E30875));
assign E30875 = (~(Vya775 | Tli675));
assign X20875 = (Joi675 & Hay775);
assign J20875 = (~(Vzu775 & Eji675));
assign H10875 = (L30875 & S30875);
assign S30875 = (~(A9i675 & Q0v775));
assign Qqr675 = (Lcz675 ? Oxh675 : hwrite_o);
assign hwrite_o = (~(Z30875 & G40875));
assign G40875 = (N40875 & U40875);
assign U40875 = (~(D7l775 & B50875));
assign B50875 = (Eh1775 | I50875);
assign I50875 = (P50875 & Rcg775);
assign P50875 = (~(F4w775 | V8p675));
assign Eh1775 = (Rfr775 & Pw9775);
assign N40875 = (~(Zx6775 & W50875));
assign W50875 = (~(Nyr775 & D60875));
assign D60875 = (~(K60875 & Zfa775));
assign K60875 = (~(K7s775 | Yaw775));
assign Nyr775 = (!Sry675);
assign Sry675 = (Nzy675 & X5p675);
assign Z30875 = (R60875 & Y60875);
assign Jqr675 = (Lcz675 ? G5i675 : F70875);
assign F70875 = (~(M70875 & T70875));
assign T70875 = (~(A80875 & H80875));
assign H80875 = (~(Q6b775 | Wxf775));
assign A80875 = (~(Yaw775 | U3g775));
assign M70875 = (~(O80875 & V80875));
assign O80875 = (~(F4w775 | Pw9775));
assign Cqr675 = (~(C90875 & J90875));
assign J90875 = (Q90875 & X90875);
assign X90875 = (~(Aft775 & Sy1l85[2]));
assign Q90875 = (Ea0875 & Oft775);
assign Ea0875 = (Vft775 | T26775);
assign T26775 = (La0875 & Sa0875);
assign Sa0875 = (Za0875 & Gb0875);
assign Gb0875 = (~(I3v775 & Nb0875));
assign Za0875 = (Ub0875 & Ufb775);
assign Ub0875 = (~(D4v775 & Bc0875));
assign La0875 = (Ic0875 & Pc0875);
assign Pc0875 = (~(F5v775 & Wc0875));
assign Ic0875 = (Yhb775 | Dd0875);
assign C90875 = (Kd0875 & Rd0875);
assign Rd0875 = (~(E52l85[1] & Ykt775));
assign Kd0875 = (~(vis_pc_o[1] & P60775));
assign Vpr675 = (~(Yd0875 & Fe0875));
assign Fe0875 = (Me0875 & Te0875);
assign Te0875 = (~(Aft775 & Sy1l85[3]));
assign Me0875 = (Af0875 & Oft775);
assign Af0875 = (Vft775 | Sx6775);
assign Sx6775 = (Hf0875 & Of0875);
assign Of0875 = (Vf0875 & Cg0875);
assign Cg0875 = (~(I3v775 & Jg0875));
assign Vf0875 = (Qg0875 & Ufb775);
assign Qg0875 = (~(D4v775 & Xg0875));
assign Hf0875 = (Eh0875 & Lh0875);
assign Lh0875 = (~(F5v775 & Sh0875));
assign Eh0875 = (Yhb775 | Zh0875);
assign Yd0875 = (Gi0875 & Ni0875);
assign Ni0875 = (~(E52l85[2] & Ykt775));
assign Gi0875 = (~(vis_pc_o[2] & P60775));
assign Opr675 = (~(Ui0875 & Bj0875));
assign Bj0875 = (Ij0875 & Pj0875);
assign Pj0875 = (~(Aft775 & Sy1l85[4]));
assign Ij0875 = (Wj0875 & Oft775);
assign Wj0875 = (Vft775 | Oh6775);
assign Oh6775 = (Dk0875 & Kk0875);
assign Kk0875 = (Rk0875 & Yk0875);
assign Yk0875 = (Zeb775 | Fl0875);
assign Rk0875 = (Ml0875 & Ufb775);
assign Ml0875 = (Bgb775 | Tl0875);
assign Dk0875 = (Am0875 & Hm0875);
assign Hm0875 = (Dhb775 | Om0875);
assign Am0875 = (Yhb775 | Vm0875);
assign Ui0875 = (Cn0875 & Jn0875);
assign Jn0875 = (~(E52l85[3] & Ykt775));
assign Cn0875 = (~(vis_pc_o[3] & P60775));
assign Hpr675 = (~(Qn0875 & Xn0875));
assign Xn0875 = (Eo0875 & Lo0875);
assign Lo0875 = (~(Aft775 & Sy1l85[5]));
assign Eo0875 = (So0875 & Oft775);
assign So0875 = (Vft775 | Mv5775);
assign Mv5775 = (Zo0875 & Gp0875);
assign Gp0875 = (Np0875 & Up0875);
assign Up0875 = (Zeb775 | Bq0875);
assign Np0875 = (Iq0875 & Ufb775);
assign Iq0875 = (Bgb775 | Pq0875);
assign Bgb775 = (!D4v775);
assign Zo0875 = (Wq0875 & Dr0875);
assign Dr0875 = (Dhb775 | Kr0875);
assign Dhb775 = (!F5v775);
assign Wq0875 = (Yhb775 | Rr0875);
assign Qn0875 = (Yr0875 & Fs0875);
assign Fs0875 = (~(E52l85[4] & Ykt775));
assign Yr0875 = (~(vis_pc_o[4] & P60775));
assign Apr675 = (~(Ms0875 & Ts0875));
assign Ts0875 = (At0875 & Ht0875);
assign Ht0875 = (~(Aft775 & Sy1l85[6]));
assign At0875 = (Ot0875 & Oft775);
assign Ot0875 = (Vft775 | Lrc775);
assign Lrc775 = (Vt0875 & Cu0875);
assign Cu0875 = (Ju0875 & Qu0875);
assign Qu0875 = (~(I3v775 & Pjt775));
assign Ju0875 = (Xu0875 & Ufb775);
assign Xu0875 = (~(D4v775 & Dkt775));
assign Vt0875 = (Ev0875 & Lv0875);
assign Lv0875 = (~(F5v775 & Lht775));
assign Ev0875 = (Nit775 | Yhb775);
assign Ms0875 = (Sv0875 & Zv0875);
assign Zv0875 = (~(E52l85[5] & Ykt775));
assign Sv0875 = (~(vis_pc_o[5] & P60775));
assign Tor675 = (~(Gw0875 & Nw0875));
assign Nw0875 = (Uw0875 & Bx0875);
assign Bx0875 = (~(Aft775 & Sy1l85[7]));
assign Uw0875 = (Ix0875 & Oft775);
assign Ix0875 = (Vft775 | N0c775);
assign N0c775 = (Px0875 & Wx0875);
assign Wx0875 = (Dy0875 & Ky0875);
assign Ky0875 = (Zeb775 | Gqz775);
assign Zeb775 = (!I3v775);
assign I3v775 = (~(Ry0875 & Yy0875));
assign Yy0875 = (~(Fz0875 & Ubm775));
assign Ry0875 = (~(Mz0875 | Tz0875));
assign Mz0875 = (A01875 & H01875);
assign A01875 = (~(O01875 | M62l85[0]));
assign Dy0875 = (V01875 & Ufb775);
assign Ufb775 = (~(C11875 & J11875));
assign J11875 = (~(Q11875 & X11875));
assign Q11875 = (~(E21875 & L21875));
assign L21875 = (S21875 & Z21875);
assign S21875 = (~(G31875 & Ubm775));
assign E21875 = (N31875 & U31875);
assign U31875 = (Tml775 | B41875);
assign Tml775 = (!Kkm775);
assign V01875 = (~(D4v775 & Qoz775));
assign D4v775 = (~(I41875 & P41875));
assign P41875 = (~(W41875 & D51875));
assign D51875 = (~(K51875 & R51875));
assign R51875 = (Y51875 & C4z675);
assign Y51875 = (~(F61875 & M61875));
assign M61875 = (~(Vxo675 & T61875));
assign T61875 = (Mwo675 | Ezo675);
assign F61875 = (~(M62l85[0] | M62l85[1]));
assign K51875 = (W1p675 & A71875);
assign A71875 = (Xza775 | Q91775);
assign Px0875 = (H71875 & O71875);
assign O71875 = (~(F5v775 & Zpz775));
assign F5v775 = (~(V71875 & C81875));
assign C81875 = (~(J81875 & M62l85[1]));
assign V71875 = (Q81875 & X81875);
assign Q81875 = (~(E91875 & Kkm775));
assign E91875 = (~(B41875 | W41875));
assign H71875 = (Epz775 | Yhb775);
assign Yhb775 = (L91875 & S91875);
assign S91875 = (Z91875 & Ga1875);
assign L91875 = (Na1875 & Ua1875);
assign Na1875 = (~(J81875 & O01875));
assign J81875 = (H01875 & M62l85[0]);
assign H01875 = (Bb1875 & W41875);
assign Bb1875 = (~(Vxo675 | X5p675));
assign Gw0875 = (Ib1875 & Pb1875);
assign Pb1875 = (~(E52l85[6] & Ykt775));
assign Ib1875 = (~(vis_pc_o[6] & P60775));
assign Mor675 = (~(Wb1875 & Dc1875));
assign Dc1875 = (Kc1875 & Rc1875);
assign Rc1875 = (~(E52l85[7] & Ykt775));
assign Kc1875 = (Yc1875 & Fd1875);
assign Fd1875 = (Vft775 | K6f775);
assign K6f775 = (Md1875 & Td1875);
assign Td1875 = (Ae1875 & He1875);
assign He1875 = (Rhb775 | Oe1875);
assign Ae1875 = (Igb775 | Ve1875);
assign Md1875 = (Cf1875 & Jf1875);
assign Jf1875 = (Gfb775 | Qf1875);
assign Cf1875 = (Khb775 | Xf1875);
assign Yc1875 = (~(Aft775 & Sy1l85[8]));
assign Wb1875 = (Eg1875 & Lg1875);
assign Lg1875 = (~(vis_pc_o[7] & P60775));
assign For675 = (~(Sg1875 & Zg1875));
assign Zg1875 = (Gh1875 & Nh1875);
assign Nh1875 = (~(Aft775 & Sy1l85[9]));
assign Gh1875 = (Uh1875 & Oft775);
assign Uh1875 = (~(Bi1875 & Aue775));
assign Aue775 = (~(Ii1875 & Pi1875));
assign Pi1875 = (Wi1875 & Dj1875);
assign Dj1875 = (~(P3v775 & Kj1875));
assign Wi1875 = (Rj1875 & Kse775);
assign Rj1875 = (~(M5v775 & Yj1875));
assign Ii1875 = (Fk1875 & Mk1875);
assign Mk1875 = (T5v775 | Oe1875);
assign Fk1875 = (~(K4v775 & Tk1875));
assign Sg1875 = (Al1875 & Hl1875);
assign Hl1875 = (~(E52l85[8] & Ykt775));
assign Al1875 = (~(vis_pc_o[8] & P60775));
assign Ynr675 = (~(Ol1875 & Vl1875));
assign Vl1875 = (Cm1875 & Jm1875);
assign Jm1875 = (~(E52l85[13] & Ykt775));
assign Cm1875 = (Qm1875 & Xm1875);
assign Xm1875 = (Vft775 | Y7e775);
assign Y7e775 = (En1875 & Ln1875);
assign Ln1875 = (Sn1875 & Zn1875);
assign Zn1875 = (~(Dkt775 & Tk1875));
assign Dkt775 = (~(Go1875 & No1875));
assign No1875 = (Uo1875 & Bp1875);
assign Bp1875 = (Ip1875 | Atm775);
assign Uo1875 = (~(Pp1875 & Wp1875));
assign Wp1875 = (~(Dq1875 & Kq1875));
assign Kq1875 = (Rq1875 & Yq1875);
assign Yq1875 = (Fr1875 & Mr1875);
assign Mr1875 = (Tr1875 & As1875);
assign As1875 = (~(Rg5775 & Mb2l85[56]));
assign Tr1875 = (~(Fh5775 & Mb2l85[48]));
assign Fr1875 = (Hs1875 & Os1875);
assign Os1875 = (~(Th5775 & Mb2l85[40]));
assign Hs1875 = (~(Hi5775 & Mb2l85[32]));
assign Rq1875 = (Vs1875 & Ct1875);
assign Ct1875 = (~(Xj5775 & Mb2l85[8]));
assign Vs1875 = (Jt1875 & Qt1875);
assign Qt1875 = (~(Vi5775 & Mb2l85[24]));
assign Jt1875 = (~(Jj5775 & Mb2l85[16]));
assign Dq1875 = (Xt1875 & Eu1875);
assign Eu1875 = (Lu1875 & Su1875);
assign Su1875 = (~(V72l85[6] & Kn5775));
assign Lu1875 = (Zu1875 & Gv1875);
assign Gv1875 = (~(Lk5775 & Mb2l85[0]));
assign Zu1875 = (~(st_calib_i[6] & Nv1875));
assign Xt1875 = (Uv1875 & Bw1875);
assign Bw1875 = (~(Iw1875 & Yg2l85[6]));
assign Uv1875 = (Pw1875 & Ww1875);
assign Ww1875 = (~(Pf2l85[6] & Wn4775));
assign Pw1875 = (~(Dx1875 & Gi2l85[6]));
assign Go1875 = (Kx1875 & Rx1875);
assign Rx1875 = (~(Yx1875 & Lvm775));
assign Kx1875 = (~(hrdata_i[6] & Fy1875));
assign Sn1875 = (Nit775 | Oe1875);
assign Nit775 = (My1875 & Ty1875);
assign Ty1875 = (Az1875 & Hz1875);
assign Hz1875 = (~(Pp1875 & Oz1875));
assign Oz1875 = (~(Vz1875 & C02875));
assign C02875 = (J02875 & Q02875);
assign Q02875 = (X02875 & E12875);
assign E12875 = (L12875 & S12875);
assign L12875 = (~(J12775 & Xqj775));
assign J12775 = (~(Z12875 | G22875));
assign Z12875 = (B32875 ? U22875 : N22875);
assign N22875 = (I32875 & P32875);
assign I32875 = (K42875 ? D42875 : W32875);
assign D42875 = (~(R42875 | Y42875));
assign Y42875 = (~(F52875 | M52875));
assign W32875 = (~(T52875 | A62875));
assign X02875 = (H62875 & O62875);
assign O62875 = (~(Rg5775 & Mb2l85[58]));
assign H62875 = (~(Fh5775 & Mb2l85[50]));
assign J02875 = (V62875 & C72875);
assign C72875 = (J72875 & Q72875);
assign Q72875 = (~(Th5775 & Mb2l85[42]));
assign J72875 = (~(Hi5775 & Mb2l85[34]));
assign V62875 = (X72875 & E82875);
assign E82875 = (~(Vi5775 & Mb2l85[26]));
assign X72875 = (~(Jj5775 & Mb2l85[18]));
assign Vz1875 = (L82875 & S82875);
assign S82875 = (Z82875 & G92875);
assign G92875 = (N92875 & U92875);
assign U92875 = (~(Xj5775 & Mb2l85[10]));
assign N92875 = (~(Lk5775 & Mb2l85[2]));
assign Z82875 = (Ba2875 & Ia2875);
assign Ia2875 = (~(st_calib_i[14] & Nv1875));
assign Ba2875 = (~(V72l85[14] & Kn5775));
assign L82875 = (Pa2875 & Wa2875);
assign Wa2875 = (~(Iw1875 & Yg2l85[14]));
assign Pa2875 = (Db2875 & Kb2875);
assign Kb2875 = (~(Pf2l85[14] & Wn4775));
assign Db2875 = (~(Dx1875 & Gi2l85[14]));
assign Az1875 = (Ip1875 | F7m775);
assign My1875 = (Rb2875 & Yb2875);
assign Yb2875 = (Fc2875 | O8m775);
assign Rb2875 = (~(hrdata_i[14] & Fy1875));
assign En1875 = (Mc2875 & Tc2875);
assign Tc2875 = (~(Pjt775 & Kj1875));
assign Pjt775 = (~(Ad2875 & Hd2875));
assign Hd2875 = (Od2875 & Vd2875);
assign Vd2875 = (Ip1875 | Rdm775);
assign Od2875 = (~(Pp1875 & Ce2875));
assign Ce2875 = (~(Je2875 & Qe2875));
assign Qe2875 = (Xe2875 & Ef2875);
assign Ef2875 = (Lf2875 & Sf2875);
assign Sf2875 = (Zf2875 & Gg2875);
assign Gg2875 = (~(Bm5775 & C92l85[0]));
assign Zf2875 = (~(Rg5775 & Mb2l85[60]));
assign Lf2875 = (Ng2875 & Ug2875);
assign Ug2875 = (~(Fh5775 & Mb2l85[52]));
assign Ng2875 = (~(Th5775 & Mb2l85[44]));
assign Xe2875 = (Bh2875 & Ih2875);
assign Ih2875 = (~(Jj5775 & Mb2l85[20]));
assign Bh2875 = (Ph2875 & Wh2875);
assign Wh2875 = (~(Hi5775 & Mb2l85[36]));
assign Ph2875 = (~(Vi5775 & Mb2l85[28]));
assign Je2875 = (Di2875 & Ki2875);
assign Ki2875 = (Ri2875 & Yi2875);
assign Yi2875 = (Fj2875 & Mj2875);
assign Mj2875 = (~(Xj5775 & Mb2l85[12]));
assign Fj2875 = (~(Lk5775 & Mb2l85[4]));
assign Ri2875 = (Tj2875 & Ak2875);
assign Ak2875 = (~(st_calib_i[22] & Nv1875));
assign Tj2875 = (~(V72l85[22] & Kn5775));
assign Di2875 = (Hk2875 & Ok2875);
assign Ok2875 = (~(Iw1875 & Yg2l85[22]));
assign Hk2875 = (Vk2875 & Cl2875);
assign Cl2875 = (~(Pf2l85[22] & Wn4775));
assign Vk2875 = (~(Dx1875 & Gi2l85[22]));
assign Ad2875 = (Jl2875 & Ql2875);
assign Ql2875 = (~(Yx1875 & Jgm775));
assign Jl2875 = (~(hrdata_i[22] & Fy1875));
assign Mc2875 = (~(Lht775 & Yj1875));
assign Lht775 = (~(Xl2875 & Em2875));
assign Em2875 = (~(Pp1875 & Lm2875));
assign Lm2875 = (~(Sm2875 & Zm2875));
assign Zm2875 = (Gn2875 & Nn2875);
assign Nn2875 = (Un2875 & Bo2875);
assign Un2875 = (Io2875 & Po2875);
assign Po2875 = (~(Nl5775 & Ha2l85[0]));
assign Io2875 = (~(Bm5775 & Ge2l85[0]));
assign Gn2875 = (Wo2875 & Dp2875);
assign Dp2875 = (Kp2875 & Rp2875);
assign Rp2875 = (~(Rg5775 & Mb2l85[62]));
assign Kp2875 = (~(Fh5775 & Mb2l85[54]));
assign Wo2875 = (Yp2875 & Fq2875);
assign Fq2875 = (~(Th5775 & Mb2l85[46]));
assign Yp2875 = (~(Hi5775 & Mb2l85[38]));
assign Sm2875 = (Mq2875 & Tq2875);
assign Tq2875 = (Ar2875 & Hr2875);
assign Hr2875 = (Or2875 & Vr2875);
assign Vr2875 = (~(Vi5775 & Mb2l85[30]));
assign Or2875 = (~(Jj5775 & Mb2l85[22]));
assign Ar2875 = (Cs2875 & Js2875);
assign Js2875 = (~(Xj5775 & Mb2l85[14]));
assign Cs2875 = (~(Lk5775 & Mb2l85[6]));
assign Mq2875 = (Qs2875 & Xs2875);
assign Xs2875 = (~(Iw1875 & Yg2l85[30]));
assign Qs2875 = (Et2875 & Lt2875);
assign Lt2875 = (~(st_calib_i[24] & Nv1875));
assign Et2875 = (~(Dx1875 & Gi2l85[30]));
assign Xl2875 = (St2875 & Zt2875);
assign Zt2875 = (~(Gu2875 & Nu2875));
assign Nu2875 = (~(Uu2875 & Bv2875));
assign Bv2875 = (Iv2875 | Lwl775);
assign Uu2875 = (~(Gpm775 & Pv2875));
assign Pv2875 = (Npm775 | Iqm775);
assign Gpm775 = (Wv2875 & Iv2875);
assign Iv2875 = (~(Dw2875 & Kw2875));
assign Dw2875 = (Fx2875 ? Yw2875 : Rw2875);
assign Wv2875 = (Mx2875 | Kll775);
assign St2875 = (~(hrdata_i[30] & Fy1875));
assign Qm1875 = (~(Aft775 & Sy1l85[14]));
assign Ol1875 = (Eg1875 & Tx2875);
assign Tx2875 = (~(vis_pc_o[13] & P60775));
assign Rnr675 = (~(Ay2875 & Hy2875));
assign Hy2875 = (Oy2875 & Vy2875);
assign Vy2875 = (~(E52l85[14] & Ykt775));
assign Oy2875 = (Cz2875 & Jz2875);
assign Jz2875 = (Vft775 | Gbf775);
assign Gbf775 = (Qz2875 & Xz2875);
assign Xz2875 = (E03875 & L03875);
assign L03875 = (~(Tk1875 & Qoz775));
assign E03875 = (Gqz775 | Qf1875);
assign Qz2875 = (S03875 & Z03875);
assign Z03875 = (~(Zpz775 & Yj1875));
assign S03875 = (Epz775 | Oe1875);
assign Cz2875 = (~(Aft775 & Sy1l85[15]));
assign Ay2875 = (Eg1875 & G13875);
assign G13875 = (~(vis_pc_o[14] & P60775));
assign Knr675 = (~(N13875 & U13875));
assign U13875 = (B23875 & I23875);
assign I23875 = (~(E52l85[15] & Ykt775));
assign B23875 = (P23875 & W23875);
assign W23875 = (Vft775 | V2e775);
assign V2e775 = (D33875 & K33875);
assign K33875 = (R33875 & Y33875);
assign Y33875 = (Ikz775 | Rhb775);
assign R33875 = (Git775 | Igb775);
assign D33875 = (F43875 & M43875);
assign M43875 = (Gfb775 | I41875);
assign F43875 = (Khb775 | T43875);
assign P23875 = (~(Aft775 & Sy1l85[16]));
assign N13875 = (Rlz775 & A53875);
assign A53875 = (~(vis_pc_o[15] & P60775));
assign Dnr675 = (~(H53875 & O53875));
assign O53875 = (V53875 & C63875);
assign C63875 = (~(E52l85[16] & Ykt775));
assign V53875 = (J63875 & Q63875);
assign Q63875 = (Vft775 | Xwd775);
assign Xwd775 = (X63875 & E73875);
assign E73875 = (L73875 & S73875);
assign S73875 = (~(M5v775 & Klz775));
assign L73875 = (~(P3v775 & Dlz775));
assign X63875 = (Z73875 & G83875);
assign G83875 = (Ikz775 | T5v775);
assign Z73875 = (~(Bkz775 & K4v775));
assign J63875 = (~(Aft775 & Sy1l85[17]));
assign H53875 = (Rlz775 & N83875);
assign N83875 = (~(vis_pc_o[16] & P60775));
assign Wmr675 = (~(U83875 & B93875));
assign B93875 = (I93875 & P93875);
assign P93875 = (~(E52l85[17] & Ykt775));
assign I93875 = (W93875 & Da3875);
assign Da3875 = (Vft775 | Urd775);
assign Urd775 = (Ka3875 & Ra3875);
assign Ra3875 = (Ya3875 & Fb3875);
assign Fb3875 = (Ikz775 | Dd0875);
assign Ya3875 = (~(Klz775 & Wc0875));
assign Ka3875 = (Mb3875 & Tb3875);
assign Tb3875 = (~(Bkz775 & Bc0875));
assign Mb3875 = (~(Nb0875 & Dlz775));
assign W93875 = (~(Aft775 & Sy1l85[18]));
assign U83875 = (Rlz775 & Ac3875);
assign Ac3875 = (~(vis_pc_o[17] & P60775));
assign Pmr675 = (~(Hc3875 & Oc3875));
assign Oc3875 = (Vc3875 & Cd3875);
assign Cd3875 = (~(E52l85[18] & Ykt775));
assign Vc3875 = (Jd3875 & Qd3875);
assign Qd3875 = (Vft775 | Ymd775);
assign Ymd775 = (Xd3875 & Ee3875);
assign Ee3875 = (Le3875 & Se3875);
assign Se3875 = (Ikz775 | Zh0875);
assign Le3875 = (~(Klz775 & Sh0875));
assign Xd3875 = (Ze3875 & Gf3875);
assign Gf3875 = (~(Bkz775 & Xg0875));
assign Ze3875 = (~(Jg0875 & Dlz775));
assign Jd3875 = (~(Aft775 & Sy1l85[19]));
assign Hc3875 = (Rlz775 & Nf3875);
assign Nf3875 = (~(vis_pc_o[18] & P60775));
assign Imr675 = (~(Uf3875 & Bg3875));
assign Bg3875 = (Ig3875 & Pg3875);
assign Pg3875 = (~(E52l85[19] & Ykt775));
assign Ig3875 = (Wg3875 & Dh3875);
assign Dh3875 = (Vft775 | Cid775);
assign Cid775 = (Kh3875 & Rh3875);
assign Rh3875 = (Yh3875 & Fi3875);
assign Fi3875 = (Ikz775 | Vm0875);
assign Yh3875 = (T43875 | Om0875);
assign Kh3875 = (Mi3875 & Ti3875);
assign Ti3875 = (Git775 | Tl0875);
assign Mi3875 = (Fl0875 | I41875);
assign Wg3875 = (~(Aft775 & Sy1l85[20]));
assign Uf3875 = (Rlz775 & Aj3875);
assign Aj3875 = (~(vis_pc_o[19] & P60775));
assign Bmr675 = (~(Hj3875 & Oj3875));
assign Oj3875 = (Vj3875 & Ck3875);
assign Ck3875 = (~(E52l85[20] & Ykt775));
assign Vj3875 = (Jk3875 & Qk3875);
assign Qk3875 = (Vft775 | Gdd775);
assign Gdd775 = (Xk3875 & El3875);
assign El3875 = (Ll3875 & Sl3875);
assign Sl3875 = (Ikz775 | Rr0875);
assign Ll3875 = (T43875 | Kr0875);
assign T43875 = (!Klz775);
assign Xk3875 = (Zl3875 & Gm3875);
assign Gm3875 = (Git775 | Pq0875);
assign Zl3875 = (I41875 | Bq0875);
assign Jk3875 = (~(Aft775 & Sy1l85[21]));
assign Hj3875 = (Rlz775 & Nm3875);
assign Nm3875 = (~(vis_pc_o[20] & P60775));
assign Ulr675 = (~(Um3875 & Bn3875));
assign Bn3875 = (In3875 & Pn3875);
assign Pn3875 = (~(Aft775 & Sy1l85[24]));
assign In3875 = (Wn3875 & Oft775);
assign Wn3875 = (Vft775 | O90775);
assign O90775 = (Do3875 & Ko3875);
assign Ko3875 = (Ro3875 & Yo3875);
assign Yo3875 = (Fp3875 | Igb775);
assign Igb775 = (Mp3875 & Tp3875);
assign Tp3875 = (~(Pp1875 & Aq3875));
assign Aq3875 = (~(Hq3875 & Oq3875));
assign Oq3875 = (Vq3875 & Cr3875);
assign Cr3875 = (~(V72l85[0] & Kn5775));
assign Vq3875 = (Jr3875 & Qr3875);
assign Qr3875 = (~(S5r675 & Pn4775));
assign Jr3875 = (~(st_calib_i[0] & Nv1875));
assign Hq3875 = (Xr3875 & Es3875);
assign Es3875 = (~(Iw1875 & Yg2l85[0]));
assign Xr3875 = (Ls3875 & Ss3875);
assign Ss3875 = (~(Pf2l85[0] & Wn4775));
assign Ls3875 = (~(Dx1875 & Gi2l85[0]));
assign Mp3875 = (Zs3875 & Gt3875);
assign Gt3875 = (Prl775 | Nt3875);
assign Prl775 = (Iqm775 ? Ut3875 : Gwm775);
assign Zs3875 = (~(hrdata_i[0] & Fy1875));
assign Ro3875 = (Bu3875 & Zht775);
assign Bu3875 = (Git775 | Rhb775);
assign Rhb775 = (Iu3875 & Pu3875);
assign Pu3875 = (~(hrdata_i[8] & Fy1875));
assign Iu3875 = (Wu3875 & Dv3875);
assign Dv3875 = (~(Pp1875 & Kv3875));
assign Kv3875 = (~(Rv3875 & Yv3875));
assign Yv3875 = (Fw3875 & Mw3875);
assign Mw3875 = (~(Pf2l85[8] & Wn4775));
assign Fw3875 = (Tw3875 & Ax3875);
assign Ax3875 = (~(st_calib_i[8] & Nv1875));
assign Tw3875 = (~(V72l85[8] & Kn5775));
assign Rv3875 = (Hx3875 & Ox3875);
assign Ox3875 = (~(Dx1875 & Gi2l85[8]));
assign Hx3875 = (~(Iw1875 & Yg2l85[8]));
assign Wu3875 = (Irl775 | Nt3875);
assign Irl775 = (Iqm775 ? Qum775 : Eam775);
assign Do3875 = (Vx3875 & Cy3875);
assign Cy3875 = (Nqz775 | Gfb775);
assign Gfb775 = (Jy3875 & Qy3875);
assign Qy3875 = (~(Pp1875 & Xy3875));
assign Xy3875 = (~(Ez3875 & Lz3875));
assign Lz3875 = (Sz3875 & Zz3875);
assign Zz3875 = (G04875 & N04875);
assign G04875 = (~(B42775 & Xqj775));
assign B42775 = (U04875 & B14875);
assign U04875 = (I14875 & K42875);
assign Sz3875 = (P14875 & W14875);
assign W14875 = (~(I1r675 & Pn4775));
assign P14875 = (~(st_calib_i[16] & Nv1875));
assign Ez3875 = (D24875 & K24875);
assign K24875 = (R24875 & Y24875);
assign Y24875 = (~(V72l85[16] & Kn5775));
assign R24875 = (~(Pf2l85[16] & Wn4775));
assign D24875 = (F34875 & M34875);
assign M34875 = (~(Dx1875 & Gi2l85[16]));
assign F34875 = (~(Iw1875 & Yg2l85[16]));
assign Jy3875 = (T34875 & A44875);
assign A44875 = (Nql775 | Nt3875);
assign Nql775 = (Iqm775 ? V8m775 : Ehm775);
assign T34875 = (~(hrdata_i[16] & Fy1875));
assign Vx3875 = (H44875 | Khb775);
assign Khb775 = (O44875 & V44875);
assign V44875 = (~(Gu2875 & C54875));
assign C54875 = (~(Cnm775 & Jnm775));
assign Jnm775 = (Gql775 | J54875);
assign Gql775 = (Kll775 ? Q54875 : Hfm775);
assign Cnm775 = (~(J54875 & Shm775));
assign J54875 = (~(Yw2875 | Zry675));
assign O44875 = (X54875 & E64875);
assign E64875 = (~(hrdata_i[24] & Fy1875));
assign X54875 = (~(Pp1875 & L64875));
assign L64875 = (~(S64875 & Z64875));
assign Z64875 = (~(Iw1875 & Yg2l85[24]));
assign S64875 = (G74875 & S12875);
assign G74875 = (~(Dx1875 & Gi2l85[24]));
assign Um3875 = (N74875 & U74875);
assign U74875 = (~(E52l85[23] & Ykt775));
assign N74875 = (~(vis_pc_o[23] & P60775));
assign Nlr675 = (~(B84875 & I84875));
assign I84875 = (P84875 & W84875);
assign W84875 = (~(Aft775 & Sy1l85[25]));
assign P84875 = (D94875 & Oft775);
assign D94875 = (Vft775 | Bmc775);
assign Bmc775 = (K94875 & R94875);
assign R94875 = (Y94875 & Fa4875);
assign Fa4875 = (~(P3v775 & Ijt775));
assign P3v775 = (~(Ma4875 & Ta4875));
assign Ta4875 = (Ab4875 & Hb4875);
assign Hb4875 = (~(Ob4875 & J9m775));
assign Ab4875 = (~(Pp1875 & Vb4875));
assign Vb4875 = (~(Cc4875 & Jc4875));
assign Jc4875 = (Qc4875 & Xc4875);
assign Xc4875 = (~(V72l85[17] & Kn5775));
assign Qc4875 = (Ed4875 & Ld4875);
assign Ld4875 = (~(K52775 & Xqj775));
assign K52775 = (Sd4875 & B14875);
assign Sd4875 = (I14875 & Zd4875);
assign Ed4875 = (~(st_calib_i[17] & Nv1875));
assign Cc4875 = (Ge4875 & Ne4875);
assign Ne4875 = (~(Iw1875 & Yg2l85[17]));
assign Ge4875 = (Ue4875 & Bf4875);
assign Bf4875 = (~(Pf2l85[17] & Wn4775));
assign Ue4875 = (~(Dx1875 & Gi2l85[17]));
assign Ma4875 = (If4875 & Pf4875);
assign Pf4875 = (Fc2875 | Ddm775);
assign If4875 = (~(hrdata_i[17] & Fy1875));
assign Y94875 = (Wf4875 & Zht775);
assign Wf4875 = (~(M5v775 & Eht775));
assign M5v775 = (~(Dg4875 & Kg4875));
assign Kg4875 = (Rg4875 & Yg4875);
assign Yg4875 = (~(Gu2875 & Fh4875));
assign Fh4875 = (~(Mh4875 & Vmm775));
assign Vmm775 = (~(Th4875 & Ai4875));
assign Th4875 = (Iqm775 ? Ofm775 : Hi4875);
assign Mh4875 = (Ai4875 | Lwl775);
assign Ai4875 = (~(Oi4875 & Vi4875));
assign Oi4875 = (Qj4875 ? Jj4875 : Cj4875);
assign Rg4875 = (Xj4875 & Ek4875);
assign Xj4875 = (Lk4875 | Sk4875);
assign Dg4875 = (Zk4875 & Gl4875);
assign Gl4875 = (~(hrdata_i[25] & Fy1875));
assign Zk4875 = (~(Nl4875 & Gi2l85[25]));
assign K94875 = (Ul4875 & Bm4875);
assign Bm4875 = (Git775 | T5v775);
assign T5v775 = (Im4875 & Pm4875);
assign Pm4875 = (Wm4875 & Dn4875);
assign Dn4875 = (~(Ob4875 & Evm775));
assign Wm4875 = (~(Pp1875 & Kn4875));
assign Kn4875 = (~(Rn4875 & Yn4875));
assign Yn4875 = (Fo4875 & Mo4875);
assign Mo4875 = (S12875 & To4875);
assign Fo4875 = (Ap4875 & Hp4875);
assign Hp4875 = (~(st_calib_i[9] & Nv1875));
assign Ap4875 = (~(V72l85[9] & Kn5775));
assign Rn4875 = (Op4875 & Vp4875);
assign Vp4875 = (~(Iw1875 & Yg2l85[9]));
assign Op4875 = (Cq4875 & Jq4875);
assign Jq4875 = (~(Pf2l85[9] & Wn4775));
assign Cq4875 = (~(Dx1875 & Gi2l85[9]));
assign Im4875 = (Qq4875 & Xq4875);
assign Xq4875 = (Fc2875 | R6m775);
assign Qq4875 = (~(hrdata_i[9] & Fy1875));
assign Ul4875 = (~(K4v775 & Wjt775));
assign K4v775 = (~(Er4875 & Lr4875));
assign Lr4875 = (Sr4875 & Zr4875);
assign Zr4875 = (Ip1875 | Gs4875);
assign Gs4875 = (!Krm775);
assign Sr4875 = (~(Pp1875 & Ns4875));
assign Ns4875 = (~(Us4875 & Bt4875));
assign Bt4875 = (It4875 & Pt4875);
assign Pt4875 = (Wt4875 & Du4875);
assign Du4875 = (~(F4r675 & Pn4775));
assign Wt4875 = (~(Zk5775 & Doh675));
assign It4875 = (Ku4875 & Ru4875);
assign Ru4875 = (~(st_calib_i[1] & Nv1875));
assign Ku4875 = (~(V72l85[1] & Kn5775));
assign Us4875 = (Yu4875 & Fv4875);
assign Fv4875 = (~(Iw1875 & Yg2l85[1]));
assign Yu4875 = (Mv4875 & Tv4875);
assign Tv4875 = (~(Pf2l85[1] & Wn4775));
assign Mv4875 = (~(Dx1875 & Gi2l85[1]));
assign Er4875 = (Aw4875 & Hw4875);
assign Hw4875 = (Fc2875 | Otm775);
assign Aw4875 = (~(hrdata_i[1] & Fy1875));
assign B84875 = (Ow4875 & Vw4875);
assign Vw4875 = (~(E52l85[24] & Ykt775));
assign Ow4875 = (~(vis_pc_o[24] & P60775));
assign Glr675 = (~(Cx4875 & Jx4875));
assign Jx4875 = (Qx4875 & Xx4875);
assign Xx4875 = (~(Aft775 & Sy1l85[26]));
assign Qx4875 = (Ey4875 & Oft775);
assign Ey4875 = (Vft775 | Wfc775);
assign Wfc775 = (Ly4875 & Sy4875);
assign Sy4875 = (Zy4875 & Gz4875);
assign Gz4875 = (~(Wjt775 & Bc0875));
assign Zy4875 = (Nz4875 & Zht775);
assign Nz4875 = (~(Eht775 & Wc0875));
assign Ly4875 = (Uz4875 & B05875);
assign B05875 = (Git775 | Dd0875);
assign Uz4875 = (~(Nb0875 & Ijt775));
assign Cx4875 = (I05875 & P05875);
assign P05875 = (~(E52l85[25] & Ykt775));
assign I05875 = (~(vis_pc_o[25] & P60775));
assign Zkr675 = (~(W05875 & D15875));
assign D15875 = (K15875 & R15875);
assign R15875 = (~(Aft775 & Sy1l85[27]));
assign K15875 = (Y15875 & Oft775);
assign Y15875 = (~(Bi1875 & Abc775));
assign Abc775 = (~(F25875 & M25875));
assign M25875 = (T25875 & A35875);
assign A35875 = (~(Wjt775 & Xg0875));
assign T25875 = (H35875 & Zht775);
assign H35875 = (~(Eht775 & Sh0875));
assign F25875 = (O35875 & V35875);
assign V35875 = (Git775 | Zh0875);
assign O35875 = (~(Jg0875 & Ijt775));
assign W05875 = (C45875 & J45875);
assign J45875 = (~(E52l85[26] & Ykt775));
assign C45875 = (~(vis_pc_o[26] & P60775));
assign Skr675 = (~(Q45875 & X45875));
assign X45875 = (E55875 & L55875);
assign L55875 = (~(Aft775 & Sy1l85[28]));
assign E55875 = (S55875 & Oft775);
assign S55875 = (Vft775 | Rz0775);
assign Rz0775 = (Z55875 & G65875);
assign G65875 = (N65875 & U65875);
assign U65875 = (Fp3875 | Tl0875);
assign N65875 = (B75875 & Zht775);
assign B75875 = (H44875 | Om0875);
assign Z55875 = (I75875 & P75875);
assign P75875 = (Git775 | Vm0875);
assign I75875 = (Fl0875 | Nqz775);
assign Q45875 = (W75875 & D85875);
assign D85875 = (~(E52l85[27] & Ykt775));
assign W75875 = (~(vis_pc_o[27] & P60775));
assign Lkr675 = (~(K85875 & R85875));
assign R85875 = (Y85875 & F95875);
assign F95875 = (~(Aft775 & Sy1l85[29]));
assign Y85875 = (M95875 & Oft775);
assign M95875 = (Vft775 | Wr0775);
assign Wr0775 = (T95875 & Aa5875);
assign Aa5875 = (Ha5875 & Oa5875);
assign Oa5875 = (Fp3875 | Pq0875);
assign Fp3875 = (!Wjt775);
assign Wjt775 = (~(Va5875 & X81875));
assign Va5875 = (~(Cb5875 & Mtl775));
assign Ha5875 = (Jb5875 & Zht775);
assign Zht775 = (~(Qb5875 & Xb5875));
assign Xb5875 = (W41875 | Nim775);
assign Nim775 = (!Ewl775);
assign Ewl775 = (~(Ec5875 & Bxm775));
assign Bxm775 = (~(Mtl775 & Lc5875));
assign Lc5875 = (Sc5875 | G31875);
assign Ec5875 = (~(Zc5875 | Jvl775));
assign Jb5875 = (H44875 | Kr0875);
assign H44875 = (!Eht775);
assign Eht775 = (~(Gd5875 & Nd5875));
assign Gd5875 = (~(Jvl775 & Z21875));
assign T95875 = (Ud5875 & Be5875);
assign Be5875 = (Git775 | Rr0875);
assign Ud5875 = (Nqz775 | Bq0875);
assign K85875 = (Ie5875 & Pe5875);
assign Pe5875 = (~(E52l85[28] & Ykt775));
assign Ie5875 = (~(vis_pc_o[28] & P60775));
assign Ekr675 = (!We5875);
assign We5875 = (hready_i ? Kf5875 : Df5875);
assign Kf5875 = (Rf5875 & Yf5875);
assign Yf5875 = (~(Fg5875 & Df5875));
assign Rf5875 = (Mg5875 & Tg5875);
assign Tg5875 = (~(H90775 & Qm2775));
assign Mg5875 = (~(Aro675 & Jl3775));
assign Df5875 = (!Spo675);
assign Xjr675 = (~(Ah5875 & Hh5875));
assign Hh5875 = (~(Oh5875 & hready_i));
assign Oh5875 = (Spo675 & Vh5875);
assign Vh5875 = (Fg5875 | W60775);
assign Ah5875 = (~(Aro675 & Ci5875));
assign Ci5875 = (P60775 | W60775);
assign Qjr675 = (L0b775 ? M1i675 : Ji5875);
assign Ji5875 = (~(Qi5875 & Xi5875));
assign Xi5875 = (Ej5875 & Lj5875);
assign Lj5875 = (J6b775 | M53775);
assign Ej5875 = (Sj5875 & Zj5875);
assign Zj5875 = (~(I2b775 & Hai675));
assign Sj5875 = (~(Cei675 & A5b775));
assign Qi5875 = (Gk5875 & Nk5875);
assign Gk5875 = (Uk5875 & Bl5875);
assign Bl5875 = (Amf775 | Q6b775);
assign Uk5875 = (Il5875 | Pl5875);
assign Jjr675 = (Wl5875 | Dm5875);
assign Dm5875 = (~(Km5875 | J5x775));
assign Wl5875 = (X5x775 ? Fzi675 : Rm5875);
assign Rm5875 = (~(Ym5875 & Fn5875));
assign Fn5875 = (On0775 | Fax775);
assign Fax775 = (~(Mn5875 | Q89775));
assign Ym5875 = (Ty2775 | K9x775);
assign Cjr675 = (Tn5875 | Ao5875);
assign Ao5875 = (~(Ho5875 | J5x775));
assign J5x775 = (Oo5875 & Qea775);
assign Qea775 = (Vo5875 & Cp5875);
assign Cp5875 = (~(Sh1775 & Miw775));
assign Vo5875 = (Olg775 | F3p675);
assign Oo5875 = (Jp5875 & Iw9775);
assign Iw9775 = (!V7g775);
assign Jp5875 = (Il5875 | Vya775);
assign Tn5875 = (X5x775 ? J0j675 : Qp5875);
assign X5x775 = (~(hready_i & Xp5875));
assign Xp5875 = (~(Eq5875 & Lq5875));
assign Lq5875 = (Sq5875 & Zq5875);
assign Zq5875 = (Gr5875 & Nr5875);
assign Nr5875 = (~(Ur5875 & Iso675));
assign Ur5875 = (~(B0z675 | C8g775));
assign Gr5875 = (Yyf775 | Sn9775);
assign Sq5875 = (Bs5875 & Is5875);
assign Is5875 = (~(Ps5875 & Zx6775));
assign Bs5875 = (H0u775 | Joi675);
assign Eq5875 = (Ws5875 & Zu9775);
assign Zu9775 = (Dt5875 & Kt5875);
assign Kt5875 = (~(Y5g775 & Clv775));
assign Dt5875 = (Rt5875 & Yt5875);
assign Yt5875 = (~(Fu5875 & Rvb775));
assign Fu5875 = (~(Mwo675 | Ezo675));
assign Rt5875 = (~(Z8a775 & D7l775));
assign Ws5875 = (Yba775 & Mu5875);
assign Mu5875 = (Zh1775 | Zfh775);
assign Yba775 = (Tu5875 & Av5875);
assign Av5875 = (Hv5875 & Ov5875);
assign Ov5875 = (Vak775 & Olg775);
assign Vak775 = (~(Vv5875 & Cm2775));
assign Hv5875 = (Cw5875 & Jw5875);
assign Jw5875 = (~(Uo9775 & Qw5875));
assign Qw5875 = (Rpi675 | Xpk775);
assign Xpk775 = (M53775 & X73775);
assign Cw5875 = (~(Xw5875 & E2u775));
assign Xw5875 = (~(Ex5875 & Lx5875));
assign Lx5875 = (~(Sx5875 | Llw775));
assign Sx5875 = (Zx5875 & Izk775);
assign Zx5875 = (~(Luu775 | C4y775));
assign Luu775 = (!Fgk775);
assign Fgk775 = (Qgi675 & Xhi675);
assign Ex5875 = (Gy5875 & Ny5875);
assign Ny5875 = (~(Gw8775 & Hk3775));
assign Gy5875 = (Ahk775 | Zqi675);
assign Tu5875 = (Uy5875 & Bz5875);
assign Bz5875 = (Iz5875 & Pz5875);
assign Pz5875 = (Wub775 | Obi675);
assign Iz5875 = (Eqk775 | H0u775);
assign H0u775 = (!Uou775);
assign Uy5875 = (~(Su9775 | Dtk775));
assign Dtk775 = (~(Jrb775 & Wz5875));
assign Wz5875 = (~(Os9775 & Xza775));
assign Jrb775 = (!D06875);
assign Su9775 = (~(K06875 & R06875));
assign R06875 = (Y06875 & Cmu775);
assign Cmu775 = (Tzt775 | Nc0775);
assign Y06875 = (~(F16875 & Nxs775));
assign F16875 = (~(Izk775 | Joi675));
assign K06875 = (M16875 & T16875);
assign T16875 = (~(A26875 & Wzr775));
assign A26875 = (~(K7s775 | Bvh675));
assign M16875 = (Wub775 | Mwo675);
assign Wub775 = (~(Fiw775 & Cg8775));
assign Qp5875 = (~(H26875 & O26875));
assign O26875 = (~(Qgi675 & Mn5875));
assign Mn5875 = (~(V26875 & C36875));
assign C36875 = (J36875 & Q36875);
assign Q36875 = (~(Q89775 & X36875));
assign X36875 = (~(Ria775 & Ia3775));
assign J36875 = (Sg9775 & Ga9775);
assign Ga9775 = (~(Rj9775 & Zfv775));
assign Rj9775 = (Sta775 & Zqi675);
assign Sg9775 = (~(Sbz775 & Ik0775));
assign V26875 = (E46875 & L46875);
assign L46875 = (~(Llw775 & Ik0775));
assign Llw775 = (Mvj775 & Tli675);
assign E46875 = (Oya775 | Lrh675);
assign H26875 = (On0775 | K9x775);
assign K9x775 = (S46875 & Ky8775);
assign S46875 = (~(Ik0775 & Sta775));
assign Ik0775 = (~(Hk3775 | Lrh675));
assign Vir675 = (L0b775 ? U2i675 : Z46875);
assign Z46875 = (~(G56875 & N56875));
assign N56875 = (U56875 & B66875);
assign B66875 = (~(I2b775 & Obi675));
assign U56875 = (I66875 & P66875);
assign P66875 = (~(W66875 & Lki675));
assign W66875 = (Jfi675 & D76875);
assign D76875 = (C89775 | Aus775);
assign I66875 = (~(D3b775 & K76875));
assign K76875 = (~(R76875 & Y76875));
assign Y76875 = (~(F86875 & F4b775));
assign F86875 = (~(Cg8775 | M86875));
assign G56875 = (Nk5875 & T86875);
assign T86875 = (Fd9775 | Q6b775);
assign Fd9775 = (!A5j675);
assign Oir675 = (Bct775 ? Iw1l85[2] : A96875);
assign Bct775 = (~(hready_i & H96875));
assign H96875 = (~(O96875 & V96875));
assign V96875 = (Ca6875 & Ja6875);
assign Ja6875 = (~(Qa6875 & E2u775));
assign Qa6875 = (~(Xa6875 & Eb6875));
assign Eb6875 = (Lb6875 & Sb6875);
assign Sb6875 = (~(Zb6875 & Bvh675));
assign Zb6875 = (Gc6875 & Nc0775);
assign Gc6875 = (~(S2u775 & Iq1775));
assign S2u775 = (~(Tli675 | Joi675));
assign Lb6875 = (Tzt775 & Qm9775);
assign Qm9775 = (~(Yfk775 & Lv8775));
assign Lv8775 = (Bni675 & Bvh675);
assign Yfk775 = (~(Hk3775 | Tli675));
assign Tzt775 = (!Hhk775);
assign Hhk775 = (Aus775 & Hk3775);
assign Xa6875 = (Nc6875 & Uc6875);
assign Uc6875 = (~(N9a775 & Bd6875));
assign Bd6875 = (Gvu775 | Hk3775);
assign Nc6875 = (C4y775 | Xhi675);
assign C4y775 = (!Bk0775);
assign Ca6875 = (~(Id6875 | Yqg775));
assign Yqg775 = (Bk0775 & Zqi675);
assign Bk0775 = (Aus775 & Tc3775);
assign Id6875 = (Pd6875 & Uo9775);
assign Uo9775 = (Nxs775 & Tc3775);
assign Pd6875 = (~(Lki675 | Xhi675));
assign O96875 = (Wd6875 & Eu9775);
assign Eu9775 = (De6875 & Ke6875);
assign Ke6875 = (~(Uou775 & Re6875));
assign Re6875 = (~(Eqk775 & Ye6875));
assign Ye6875 = (Orv775 | Ff6875);
assign Orv775 = (Nh9775 | Xhi675);
assign Nh9775 = (!U3u775);
assign Eqk775 = (!W4u775);
assign W4u775 = (Lki675 & X73775);
assign Uou775 = (Nxs775 & Hk3775);
assign De6875 = (~(D06875 | Sbz775));
assign Sbz775 = (Mvj775 & Zqi675);
assign Mvj775 = (Aus775 & Ye0775);
assign D06875 = (~(Dj9775 | Wnb775));
assign Wd6875 = (Mf6875 & Fca775);
assign Fca775 = (B0z675 | Veg775);
assign Mf6875 = (~(Dba775 & D1z675));
assign A96875 = (~(Tf6875 & Ag6875));
assign Ag6875 = (Hg6875 & Og6875);
assign Og6875 = (~(Vzu775 & Lki675));
assign Vzu775 = (~(Vg6875 | Vya775));
assign Vg6875 = (Zqi675 ? Hk3775 : Ch6875);
assign Ch6875 = (Ye0775 | Rpi675);
assign Hg6875 = (~(C0v775 & Cei675));
assign C0v775 = (Eew775 & Jh6875);
assign Jh6875 = (~(Qh6875 & F6u775));
assign F6u775 = (!Ous775);
assign Qh6875 = (Joi675 ? Ei6875 : Xh6875);
assign Ei6875 = (~(Ria775 & Eji675));
assign Xh6875 = (Ef3775 ? Rpi675 : Zqi675);
assign Tf6875 = (Ict775 & Li6875);
assign Li6875 = (~(Hai675 & Q0v775));
assign Q0v775 = (Rdt775 | Si6875);
assign Si6875 = (Ddt775 & Xt2775);
assign Ict775 = (Zi6875 & Gj6875);
assign Gj6875 = (Nj6875 & Uj6875);
assign Uj6875 = (~(X5p675 & Bk6875));
assign Bk6875 = (Zry675 | Obi675);
assign Nj6875 = (Ik6875 & Dj9775);
assign Dj9775 = (!N3g775);
assign N3g775 = (Lrh675 & Cg8775);
assign Ik6875 = (~(Ria775 & Pk6875));
assign Pk6875 = (X73775 | Ye0775);
assign Ye0775 = (!Joi675);
assign X73775 = (!Eji675);
assign Zi6875 = (L30875 & Wk6875);
assign Wk6875 = (~(Joi675 & Hay775));
assign L30875 = (Dl6875 & Kl6875);
assign Kl6875 = (~(Rdt775 & Rl6875));
assign Rl6875 = (~(Tc3775 & Ply775));
assign Ply775 = (Gvu775 | M53775);
assign Gvu775 = (!Izk775);
assign Rdt775 = (Yl6875 & Fm6875);
assign Fm6875 = (Mm6875 & Ef3775);
assign Mm6875 = (~(Joi675 | Zqi675));
assign Dl6875 = (Tm6875 & Eot775);
assign Eot775 = (~(Yl6875 & Ria775));
assign Yl6875 = (~(Hk3775 | Vya775));
assign Tm6875 = (~(An6875 & Ora775));
assign Ora775 = (Fm0775 & Dr1775);
assign Dr1775 = (!A9i675);
assign Fm0775 = (!T7i675);
assign An6875 = (Obi675 & Ddt775);
assign Hir675 = (L0b775 ? Wyh675 : Hn6875);
assign L0b775 = (~(hready_i & On6875));
assign On6875 = (~(Vn6875 & Co6875));
assign Co6875 = (Jo6875 & Qo6875);
assign Qo6875 = (Xo6875 & Ep6875);
assign Ep6875 = (~(Lp6875 & U2a775));
assign U2a775 = (Sp6875 & Sta775);
assign Sp6875 = (~(Lrh675 | Zqi675));
assign Lp6875 = (Zp6875 & E2u775);
assign Zp6875 = (Rpi675 | D6t775);
assign D6t775 = (Tli675 & Ia3775);
assign Xo6875 = (Y3w775 & Vl9775);
assign Vl9775 = (~(Gq6875 & Zsb775));
assign Zsb775 = (~(Fkg775 | N0p675));
assign Gq6875 = (~(Rba775 | U50775));
assign Y3w775 = (B2b775 | Zry675);
assign B2b775 = (!Unv775);
assign Jo6875 = (Nq6875 & Uq6875);
assign Uq6875 = (~(Y5g775 & Br6875));
assign Br6875 = (Clv775 | Lrh675);
assign Clv775 = (!O6a775);
assign Y5g775 = (~(Ln9775 | Fkg775));
assign Nq6875 = (Ir6875 & Pr6875);
assign Pr6875 = (~(Jos775 & Miw775));
assign Jos775 = (~(Q91775 | Ezo675));
assign Ir6875 = (~(Wk0775 & Wr6875));
assign Wr6875 = (T1s775 | D7l775);
assign D7l775 = (Zck775 & O4p675);
assign Wk0775 = (~(Vya775 | Bvh675));
assign Vn6875 = (Ds6875 & Ks6875);
assign Ks6875 = (Rs6875 & Ys6875);
assign Ys6875 = (Zyx775 | Xt2775);
assign Xt2775 = (!Obi675);
assign Zyx775 = (~(Ft6875 & Fiw775));
assign Fiw775 = (Mt6875 & Tt6875);
assign Tt6875 = (~(Rpi675 | Ezo675));
assign Mt6875 = (Jf9775 & Hay775);
assign Ft6875 = (~(Vya775 | Mwo675));
assign Rs6875 = (Au6875 & Hu6875);
assign Hu6875 = (~(Ou6875 & E5z675));
assign Ou6875 = (~(Vu6875 & Cv6875));
assign Cv6875 = (Il5875 | Jv6875);
assign Vu6875 = (~(Gw8775 & Ib9775));
assign Ib9775 = (~(Jqx775 | Hk3775));
assign Gw8775 = (N9a775 & Tc3775);
assign Au6875 = (~(Qv6875 & Tc3775));
assign Tc3775 = (!Tli675);
assign Qv6875 = (~(Xv6875 & Ew6875));
assign Ew6875 = (~(Lw6875 & Sw6875));
assign Sw6875 = (Zw6875 & U3u775);
assign U3u775 = (Eji675 & Ia3775);
assign Zw6875 = (~(Si0775 | Cei675));
assign Si0775 = (M53775 | Ef3775);
assign M53775 = (!Xhi675);
assign Lw6875 = (~(Lyj775 | Ky8775));
assign Ky8775 = (~(Gx6875 & Ous775));
assign Ous775 = (Joi675 & Rpi675);
assign Gx6875 = (Nxs775 & E5z675);
assign Nxs775 = (Zqi675 & Bvh675);
assign Lyj775 = (!Ff6875);
assign Ff6875 = (Qgi675 & On0775);
assign Xv6875 = (~(Nx6875 & Ux6875));
assign Ux6875 = (Q89775 & Izk775);
assign Izk775 = (Lki675 & Eji675);
assign Q89775 = (C89775 & Zfv775);
assign Nx6875 = (Mpw775 & Ria775);
assign Ria775 = (~(Nc0775 | Ef3775));
assign Mpw775 = (By6875 & Ilk775);
assign By6875 = (~(Ty2775 | Xhi675));
assign Ds6875 = (Y60875 & Iy6875);
assign Iy6875 = (~(Os9775 & Zck775));
assign Y60875 = (Olg775 & Py6875);
assign Py6875 = (~(Ons775 & Rcg775));
assign Hn6875 = (~(Wy6875 & Dz6875));
assign Dz6875 = (Kz6875 & Rz6875);
assign Rz6875 = (~(Obi675 & A5b775));
assign A5b775 = (~(Whv775 & Yz6875));
assign Yz6875 = (Ahk775 | Ia3775);
assign Ia3775 = (!Lki675);
assign Whv775 = (!Aus775);
assign Aus775 = (Bvh675 & Ef3775);
assign Ef3775 = (!Bni675);
assign Kz6875 = (F07875 & M07875);
assign M07875 = (~(I2b775 & T7i675));
assign I2b775 = (~(Ahk775 | Lki675));
assign Ahk775 = (!C89775);
assign C89775 = (Joi675 & Bvh675);
assign F07875 = (~(D3b775 & T07875));
assign T07875 = (~(A17875 & H17875));
assign H17875 = (O17875 & V17875);
assign V17875 = (C27875 | Qos775);
assign Qos775 = (!R76875);
assign R76875 = (C27875 | J0j675);
assign O17875 = (~(M86875 & Y3b775));
assign A17875 = (J27875 & Q27875);
assign Q27875 = (T4b775 | F4b775);
assign J27875 = (B49775 | N1j675);
assign Wy6875 = (X27875 & Nk5875);
assign Nk5875 = (E37875 & O5b775);
assign O5b775 = (Ct9775 & Lvf775);
assign Lvf775 = (Eta775 | K1z675);
assign Ct9775 = (Fkg775 | K1z675);
assign Fkg775 = (!My9775);
assign E37875 = (~(Unv775 | Jf9775));
assign X27875 = (L37875 & S37875);
assign S37875 = (J6b775 | On0775);
assign On0775 = (!Jfi675);
assign J6b775 = (!Sta775);
assign Sta775 = (N9a775 & Bni675);
assign N9a775 = (~(Cm2775 | Joi675));
assign L37875 = (Bx8775 | Q6b775);
assign Air675 = (~(Z37875 & G47875));
assign G47875 = (N47875 & U47875);
assign U47875 = (~(E52l85[22] & Ykt775));
assign N47875 = (B57875 & I57875);
assign I57875 = (Vft775 | Qfg775);
assign Qfg775 = (P57875 & W57875);
assign W57875 = (D67875 & K67875);
assign K67875 = (Ikz775 | Epz775);
assign Ikz775 = (X81875 & R67875);
assign D67875 = (~(Klz775 & Zpz775));
assign Klz775 = (Y67875 | Cb5875);
assign P57875 = (F77875 & M77875);
assign M77875 = (~(Bkz775 & Qoz775));
assign Bkz775 = (!Git775);
assign F77875 = (Gqz775 | I41875);
assign B57875 = (~(Aft775 & Sy1l85[23]));
assign Z37875 = (Rlz775 & T77875);
assign T77875 = (~(vis_pc_o[22] & P60775));
assign Rlz775 = (Oft775 & A87875);
assign A87875 = (J3e775 | Vft775);
assign J3e775 = (~(H87875 & Qb5875));
assign Qb5875 = (O87875 & C11875);
assign O87875 = (~(V87875 & C97875));
assign C97875 = (J97875 & X11875);
assign J97875 = (~(Q97875 & T5a775));
assign Q97875 = (~(Cm2775 | U50775));
assign V87875 = (W41875 & X97875);
assign X97875 = (~(F3p675 & Kny675));
assign H87875 = (Ea7875 & Git775);
assign Git775 = (~(Fz0875 & Mtl775));
assign Ea7875 = (~(La7875 & Z21875));
assign La7875 = (~(Sa7875 & Uwm775));
assign Sa7875 = (~(Sc5875 | Zc5875));
assign Zc5875 = (!Swl775);
assign Thr675 = (~(Za7875 & Gb7875));
assign Gb7875 = (Nb7875 & Ub7875);
assign Ub7875 = (~(E52l85[9] & Ykt775));
assign Nb7875 = (Bc7875 & Ic7875);
assign Ic7875 = (Vft775 | Wre775);
assign Wre775 = (Pc7875 & Wc7875);
assign Wc7875 = (Dd7875 & Kd7875);
assign Kd7875 = (~(Bc0875 & Tk1875));
assign Bc0875 = (~(Rd7875 & Yd7875));
assign Yd7875 = (Fe7875 & Me7875);
assign Me7875 = (Ip1875 | Te7875);
assign Te7875 = (!Npm775);
assign Npm775 = (~(Af7875 & Hf7875));
assign Hf7875 = (Of7875 & Vf7875);
assign Vf7875 = (Cg7875 | Ify675);
assign Of7875 = (Jg7875 | Dgy675);
assign Af7875 = (Qg7875 & Xg7875);
assign Xg7875 = (~(Eh7875 & Lh7875));
assign Qg7875 = (Sh7875 | Bfy675);
assign Fe7875 = (~(Pp1875 & Zh7875));
assign Zh7875 = (~(Gi7875 & Ni7875));
assign Ni7875 = (Ui7875 & Bj7875);
assign Bj7875 = (Ij7875 & Pj7875);
assign Pj7875 = (~(Pn4775 & L8h775));
assign L8h775 = (S2r675 | st_calib_i[25]);
assign Pn4775 = (~(Wj7875 | Hr3775));
assign Ij7875 = (~(Fap675 & Zk5775));
assign Ui7875 = (Dk7875 & Kk7875);
assign Kk7875 = (~(st_calib_i[2] & Nv1875));
assign Dk7875 = (~(V72l85[2] & Kn5775));
assign Gi7875 = (Rk7875 & Yk7875);
assign Yk7875 = (~(Iw1875 & Yg2l85[2]));
assign Rk7875 = (Fl7875 & Ml7875);
assign Ml7875 = (~(Pf2l85[2] & Wn4775));
assign Fl7875 = (~(Dx1875 & Gi2l85[2]));
assign Rd7875 = (Tl7875 & Am7875);
assign Am7875 = (Fc2875 | Atm775);
assign Atm775 = (Hm7875 & Om7875);
assign Om7875 = (Vm7875 & Cn7875);
assign Cn7875 = (~(Eh7875 & Jn7875));
assign Vm7875 = (Cg7875 | Gey675);
assign Hm7875 = (Qn7875 & Xn7875);
assign Xn7875 = (Sh7875 | Zdy675);
assign Qn7875 = (Jg7875 | Ney675);
assign Tl7875 = (~(hrdata_i[2] & Fy1875));
assign Dd7875 = (Dd0875 | Oe1875);
assign Dd0875 = (Eo7875 & Lo7875);
assign Lo7875 = (So7875 & Zo7875);
assign Zo7875 = (~(Ob4875 & Lvm775));
assign Lvm775 = (~(Gp7875 & Np7875));
assign Np7875 = (Up7875 & Bq7875);
assign Bq7875 = (Cg7875 | Nly675);
assign Up7875 = (Sh7875 | Gly675);
assign Gp7875 = (Iq7875 & Pq7875);
assign Pq7875 = (~(Eh7875 & Wq7875));
assign Iq7875 = (Jg7875 | Uly675);
assign So7875 = (~(Pp1875 & Dr7875));
assign Dr7875 = (~(Kr7875 & Rr7875));
assign Rr7875 = (Yr7875 & Fs7875);
assign Fs7875 = (~(Pf2l85[10] & Wn4775));
assign Yr7875 = (Ms7875 & Ts7875);
assign Ts7875 = (~(st_calib_i[10] & Nv1875));
assign Ms7875 = (~(V72l85[10] & Kn5775));
assign Kr7875 = (At7875 & Ht7875);
assign Ht7875 = (~(Dx1875 & Gi2l85[10]));
assign At7875 = (~(Iw1875 & Yg2l85[10]));
assign Eo7875 = (Ot7875 & Vt7875);
assign Vt7875 = (Fc2875 | F7m775);
assign F7m775 = (Cu7875 & Ju7875);
assign Ju7875 = (Qu7875 & Xu7875);
assign Xu7875 = (~(Eh7875 & Ev7875));
assign Qu7875 = (Cg7875 | Lky675);
assign Cu7875 = (Lv7875 & Sv7875);
assign Sv7875 = (Sh7875 | Eky675);
assign Lv7875 = (Jg7875 | Sky675);
assign Ot7875 = (~(hrdata_i[10] & Fy1875));
assign Pc7875 = (Zv7875 & Gw7875);
assign Gw7875 = (~(Nb0875 & Kj1875));
assign Nb0875 = (~(Nw7875 & Uw7875));
assign Uw7875 = (Bx7875 & Ix7875);
assign Ix7875 = (Ip1875 | O8m775);
assign O8m775 = (Px7875 & Wx7875);
assign Wx7875 = (Dy7875 & Ky7875);
assign Ky7875 = (~(Eh7875 & Ry7875));
assign Dy7875 = (Sh7875 | Viy675);
assign Px7875 = (Yy7875 & Fz7875);
assign Fz7875 = (Cg7875 | Jjy675);
assign Yy7875 = (Jg7875 | Qjy675);
assign Bx7875 = (~(Pp1875 & Mz7875));
assign Mz7875 = (~(Tz7875 & A08875));
assign A08875 = (H08875 & Bo2875);
assign Bo2875 = (S12875 & N04875);
assign H08875 = (O08875 & V08875);
assign V08875 = (~(st_calib_i[18] & Nv1875));
assign O08875 = (~(V72l85[18] & Kn5775));
assign Tz7875 = (C18875 & J18875);
assign J18875 = (~(Iw1875 & Yg2l85[18]));
assign C18875 = (Q18875 & X18875);
assign X18875 = (~(Pf2l85[18] & Wn4775));
assign Q18875 = (~(Dx1875 & Gi2l85[18]));
assign Nw7875 = (E28875 & L28875);
assign L28875 = (Fc2875 | Rdm775);
assign Rdm775 = (S28875 & Z28875);
assign Z28875 = (G38875 & N38875);
assign N38875 = (~(Eh7875 & U38875));
assign G38875 = (Cg7875 | Aiy675);
assign S28875 = (B48875 & I48875);
assign I48875 = (Sh7875 | Thy675);
assign B48875 = (Jg7875 | Hiy675);
assign E28875 = (~(hrdata_i[18] & Fy1875));
assign Zv7875 = (~(Wc0875 & Yj1875));
assign Wc0875 = (~(P48875 & W48875));
assign W48875 = (~(Pp1875 & D58875));
assign D58875 = (~(K58875 & R58875));
assign R58875 = (~(Iw1875 & Yg2l85[26]));
assign K58875 = (Y58875 & F68875);
assign F68875 = (~(E7r675 & Xqj775));
assign Y58875 = (~(Dx1875 & Gi2l85[26]));
assign P48875 = (M68875 & T68875);
assign T68875 = (~(Gu2875 & A78875));
assign A78875 = (~(H78875 & Qnm775));
assign Qnm775 = (~(O78875 & V78875));
assign O78875 = (Iqm775 ? Jgm775 : Mx2875);
assign Jgm775 = (~(C88875 & J88875));
assign J88875 = (Q88875 & X88875);
assign X88875 = (~(Eh7875 & E98875));
assign Q88875 = (Sh7875 | Rgy675);
assign C88875 = (L98875 & S98875);
assign S98875 = (Cg7875 | Ygy675);
assign L98875 = (Jg7875 | Fhy675);
assign Mx2875 = (~(Z98875 & Ga8875));
assign Ga8875 = (Na8875 & Ua8875);
assign Ua8875 = (~(Eh7875 & Bb8875));
assign Na8875 = (Sh7875 | Bmy675);
assign Z98875 = (Ib8875 & Pb8875);
assign Pb8875 = (Cg7875 | Pfy675);
assign Ib8875 = (Jg7875 | Wfy675);
assign H78875 = (V78875 | Lwl775);
assign V78875 = (~(Wb8875 & Vi4875));
assign Wb8875 = (Fx2875 ? Jj4875 : Cj4875);
assign M68875 = (~(hrdata_i[26] & Fy1875));
assign Bc7875 = (~(Aft775 & Sy1l85[10]));
assign Za7875 = (Eg1875 & Dc8875);
assign Dc8875 = (~(vis_pc_o[9] & P60775));
assign Mhr675 = (~(Kc8875 & Rc8875));
assign Rc8875 = (Yc8875 & Fd8875);
assign Fd8875 = (~(E52l85[10] & Ykt775));
assign Yc8875 = (Md8875 & Td8875);
assign Td8875 = (Vft775 | Lpe775);
assign Lpe775 = (Ae8875 & He8875);
assign He8875 = (Oe8875 & Ve8875);
assign Ve8875 = (~(Xg0875 & Tk1875));
assign Tk1875 = (!Ve1875);
assign Xg0875 = (~(Cf8875 & Jf8875));
assign Jf8875 = (Qf8875 & Xf8875);
assign Xf8875 = (Fc2875 | Xum775);
assign Qf8875 = (~(Pp1875 & Eg8875));
assign Eg8875 = (~(Lg8875 & Sg8875));
assign Sg8875 = (Zg8875 & Gh8875);
assign Gh8875 = (~(V72l85[3] & Kn5775));
assign Zg8875 = (Nh8875 & To4875);
assign To4875 = (~(Uh8875 & Bi8875));
assign Uh8875 = (~(Ii8875 | Aar675));
assign Nh8875 = (~(st_calib_i[3] & Nv1875));
assign Lg8875 = (Pi8875 & Wi8875);
assign Wi8875 = (~(Iw1875 & Yg2l85[3]));
assign Pi8875 = (Dj8875 & Kj8875);
assign Kj8875 = (~(Pf2l85[3] & Wn4775));
assign Dj8875 = (~(Dx1875 & Gi2l85[3]));
assign Cf8875 = (Rj8875 & Yj8875);
assign Yj8875 = (Ip1875 | Dll775);
assign Rj8875 = (~(hrdata_i[3] & Fy1875));
assign Oe8875 = (Zh0875 | Oe1875);
assign Zh0875 = (Fk8875 & Mk8875);
assign Mk8875 = (Tk8875 & Al8875);
assign Al8875 = (Ip1875 | Lam775);
assign Tk8875 = (~(Pp1875 & Hl8875));
assign Hl8875 = (~(Ol8875 & Vl8875));
assign Vl8875 = (Cm8875 & Jm8875);
assign Jm8875 = (~(Pf2l85[11] & Wn4775));
assign Cm8875 = (Qm8875 & Xm8875);
assign Xm8875 = (~(st_calib_i[11] & Nv1875));
assign Qm8875 = (~(V72l85[11] & Kn5775));
assign Ol8875 = (En8875 & Ln8875);
assign Ln8875 = (~(Dx1875 & Gi2l85[11]));
assign En8875 = (~(Iw1875 & Yg2l85[11]));
assign Fk8875 = (Sn8875 & Zn8875);
assign Zn8875 = (~(Yx1875 & C9m775));
assign Sn8875 = (~(hrdata_i[11] & Fy1875));
assign Ae8875 = (Go8875 & No8875);
assign No8875 = (~(Jg0875 & Kj1875));
assign Jg0875 = (~(Uo8875 & Bp8875));
assign Bp8875 = (Ip8875 & Pp8875);
assign Pp8875 = (Fc2875 | Vfm775);
assign Ip8875 = (~(Pp1875 & Wp8875));
assign Wp8875 = (~(Dq8875 & Kq8875));
assign Kq8875 = (Rq8875 & Yq8875);
assign Yq8875 = (~(V72l85[19] & Kn5775));
assign Rq8875 = (Fr8875 & S12875);
assign Fr8875 = (~(st_calib_i[19] & Nv1875));
assign Dq8875 = (Mr8875 & Tr8875);
assign Tr8875 = (~(Iw1875 & Yg2l85[19]));
assign Mr8875 = (As8875 & Hs8875);
assign Hs8875 = (~(Pf2l85[19] & Wn4775));
assign As8875 = (~(Dx1875 & Gi2l85[19]));
assign Uo8875 = (Os8875 & Vs8875);
assign Vs8875 = (~(Ob4875 & Lhm775));
assign Os8875 = (~(hrdata_i[19] & Fy1875));
assign Go8875 = (~(Sh0875 & Yj1875));
assign Sh0875 = (~(Ct8875 & Jt8875));
assign Jt8875 = (Qt8875 & Xt8875);
assign Xt8875 = (~(Nl4875 & Gi2l85[27]));
assign Qt8875 = (Eu8875 & Ek4875);
assign Eu8875 = (~(hrdata_i[27] & Fy1875));
assign Ct8875 = (Lu8875 & Su8875);
assign Su8875 = (~(Gu2875 & Zu8875));
assign Zu8875 = (~(Gv8875 & Bqm775));
assign Bqm775 = (Nv8875 | Uv8875);
assign Nv8875 = (Kll775 ? Wkl775 : Bw8875);
assign Gv8875 = (~(Uv8875 & Shm775));
assign Uv8875 = (Iw8875 & Vi4875);
assign Vi4875 = (Ezo675 & Rw2875);
assign Iw8875 = (Jg7875 ? Jj4875 : Cj4875);
assign Lu8875 = (Lk4875 | Pw8875);
assign Md8875 = (~(Aft775 & Sy1l85[11]));
assign Kc8875 = (Eg1875 & Ww8875);
assign Ww8875 = (~(vis_pc_o[10] & P60775));
assign Fhr675 = (~(Dx8875 & Kx8875));
assign Kx8875 = (Rx8875 & Yx8875);
assign Yx8875 = (~(E52l85[11] & Ykt775));
assign Rx8875 = (Fy8875 & My8875);
assign My8875 = (Vft775 | Zie775);
assign Zie775 = (Ty8875 & Az8875);
assign Az8875 = (Hz8875 & Oz8875);
assign Oz8875 = (Tl0875 | Ve1875);
assign Tl0875 = (Vz8875 & C09875);
assign C09875 = (J09875 & Q09875);
assign Q09875 = (Fc2875 | Qum775);
assign Qum775 = (X09875 & E19875);
assign E19875 = (L19875 & S19875);
assign S19875 = (Cg7875 | Sdy675);
assign L19875 = (Jg7875 | Zdy675);
assign X09875 = (Z19875 & G29875);
assign G29875 = (N29875 | Nly675);
assign Z19875 = (Sh7875 | Uly675);
assign J09875 = (~(Pp1875 & U29875));
assign U29875 = (~(B39875 & I39875));
assign I39875 = (P39875 & W39875);
assign W39875 = (~(V72l85[4] & Kn5775));
assign P39875 = (D49875 & K49875);
assign K49875 = (~(Nbp675 & Zk5775));
assign Zk5775 = (R49875 & Y49875);
assign R49875 = (~(F59875 | Aar675));
assign D49875 = (~(st_calib_i[4] & Nv1875));
assign B39875 = (M59875 & T59875);
assign T59875 = (~(Iw1875 & Yg2l85[4]));
assign M59875 = (A69875 & H69875);
assign H69875 = (~(Pf2l85[4] & Wn4775));
assign A69875 = (~(Dx1875 & Gi2l85[4]));
assign Vz8875 = (O69875 & V69875);
assign V69875 = (Ip1875 | Gwm775);
assign Gwm775 = (C79875 & J79875);
assign J79875 = (Q79875 & X79875);
assign X79875 = (~(Eh7875 & E89875));
assign Q79875 = (Sh7875 | Ney675);
assign C79875 = (L89875 & S89875);
assign S89875 = (Cg7875 | Uey675);
assign L89875 = (Jg7875 | Bfy675);
assign O69875 = (~(hrdata_i[4] & Fy1875));
assign Hz8875 = (Vm0875 | Oe1875);
assign Vm0875 = (Z89875 & G99875);
assign G99875 = (N99875 & U99875);
assign U99875 = (Fc2875 | V8m775);
assign V8m775 = (Ba9875 & Ia9875);
assign Ia9875 = (Pa9875 & Wa9875);
assign Wa9875 = (Jg7875 | Eky675);
assign Pa9875 = (N29875 | Jjy675);
assign Ba9875 = (Db9875 & Kb9875);
assign Kb9875 = (Sh7875 | Qjy675);
assign Db9875 = (Cg7875 | Xjy675);
assign N99875 = (~(Pp1875 & Rb9875));
assign Rb9875 = (~(Yb9875 & Fc9875));
assign Fc9875 = (Mc9875 & Tc9875);
assign Tc9875 = (~(V72l85[12] & Kn5775));
assign Mc9875 = (Ad9875 & Hd9875);
assign Hd9875 = (~(Ju1775 & Xqj775));
assign Ju1775 = (Od9875 & Vpj775);
assign Od9875 = (Vd9875 | Cep675);
assign Vd9875 = (B32875 ? U22875 : Ce9875);
assign Ce9875 = (~(P32875 & Je9875));
assign Je9875 = (~(Qe9875 & Xe9875));
assign Qe9875 = (K42875 ? Lf9875 : Ef9875);
assign Lf9875 = (Gg9875 ? Zf9875 : Sf9875);
assign Zf9875 = (M52875 ? Ug9875 : Ng9875);
assign Ug9875 = (Ph9875 ? Ih9875 : Bh9875);
assign Ng9875 = (Ki9875 ? Di9875 : Wh9875);
assign Sf9875 = (Fj9875 ? Yi9875 : Ri9875);
assign Yi9875 = (Ak9875 ? Tj9875 : Mj9875);
assign Ri9875 = (Vk9875 ? Ok9875 : Hk9875);
assign Ef9875 = (Ql9875 ? Jl9875 : Cl9875);
assign Jl9875 = (Lm9875 ? Em9875 : Xl9875);
assign Em9875 = (Gn9875 ? Zm9875 : Sm9875);
assign Xl9875 = (Bo9875 ? Un9875 : Nn9875);
assign Cl9875 = (Wo9875 ? Po9875 : Io9875);
assign Po9875 = (Rp9875 ? Kp9875 : Dp9875);
assign Io9875 = (Mq9875 ? Fq9875 : Yp9875);
assign Ad9875 = (~(st_calib_i[12] & Nv1875));
assign Yb9875 = (Tq9875 & Ar9875);
assign Ar9875 = (~(Iw1875 & Yg2l85[12]));
assign Tq9875 = (Hr9875 & Or9875);
assign Or9875 = (~(Pf2l85[12] & Wn4775));
assign Hr9875 = (~(Dx1875 & Gi2l85[12]));
assign Z89875 = (Vr9875 & Cs9875);
assign Cs9875 = (Ip1875 | Eam775);
assign Eam775 = (Js9875 & Qs9875);
assign Qs9875 = (Xs9875 & Et9875);
assign Et9875 = (Jg7875 | Gly675);
assign Xs9875 = (N29875 | Lky675);
assign Js9875 = (Lt9875 & St9875);
assign St9875 = (Sh7875 | Sky675);
assign Lt9875 = (Cg7875 | Zky675);
assign Vr9875 = (~(hrdata_i[12] & Fy1875));
assign Ty8875 = (Zt9875 & Gu9875);
assign Gu9875 = (Fl0875 | Qf1875);
assign Fl0875 = (Nu9875 & Uu9875);
assign Uu9875 = (Bv9875 & Iv9875);
assign Iv9875 = (Ip1875 | Ehm775);
assign Ehm775 = (Pv9875 & Wv9875);
assign Wv9875 = (Dw9875 & Kw9875);
assign Kw9875 = (N29875 | Aiy675);
assign Dw9875 = (Sh7875 | Hiy675);
assign Pv9875 = (Rw9875 & Yw9875);
assign Yw9875 = (Cg7875 | Oiy675);
assign Rw9875 = (Jg7875 | Viy675);
assign Bv9875 = (~(Pp1875 & Fx9875));
assign Fx9875 = (~(Mx9875 & Tx9875));
assign Tx9875 = (Ay9875 & Hy9875);
assign Hy9875 = (~(Pf2l85[20] & Wn4775));
assign Ay9875 = (Oy9875 & Vy9875);
assign Vy9875 = (~(st_calib_i[20] & Nv1875));
assign Oy9875 = (~(V72l85[20] & Kn5775));
assign Mx9875 = (Cz9875 & Jz9875);
assign Jz9875 = (~(Dx1875 & Gi2l85[20]));
assign Cz9875 = (~(Iw1875 & Yg2l85[20]));
assign Nu9875 = (Qz9875 & Xz9875);
assign Xz9875 = (Fc2875 | Hfm775);
assign Hfm775 = (E0a875 & L0a875);
assign L0a875 = (S0a875 & Z0a875);
assign Z0a875 = (N29875 | Ygy675);
assign S0a875 = (Jg7875 | Thy675);
assign E0a875 = (G1a875 & N1a875);
assign N1a875 = (Cg7875 | Mhy675);
assign G1a875 = (Sh7875 | Fhy675);
assign Fc2875 = (!Yx1875);
assign Qz9875 = (~(hrdata_i[20] & Fy1875));
assign Zt9875 = (Om0875 | Xf1875);
assign Om0875 = (U1a875 & B2a875);
assign B2a875 = (I2a875 & Ek4875);
assign I2a875 = (~(Pp1875 & P2a875));
assign P2a875 = (~(W2a875 & D3a875));
assign D3a875 = (~(Iw1875 & Yg2l85[28]));
assign W2a875 = (K3a875 & R3a875);
assign R3a875 = (~(Ifp675 & Xqj775));
assign K3a875 = (~(Dx1875 & Gi2l85[28]));
assign U1a875 = (Y3a875 & F4a875);
assign F4a875 = (~(Gu2875 & M4a875));
assign M4a875 = (~(T4a875 & Xnm775));
assign Xnm775 = (A5a875 | H5a875);
assign A5a875 = (Kll775 ? Ut3875 : Q54875);
assign Ut3875 = (O5a875 & V5a875);
assign V5a875 = (C6a875 & J6a875);
assign J6a875 = (~(Eh7875 & Q6a875));
assign C6a875 = (Sh7875 | Dgy675);
assign O5a875 = (X6a875 & E7a875);
assign E7a875 = (Cg7875 | Cjy675);
assign X6a875 = (Jg7875 | Bmy675);
assign Q54875 = (L7a875 & S7a875);
assign S7a875 = (Z7a875 & G8a875);
assign G8a875 = (Sh7875 | Wfy675);
assign Z7a875 = (Jg7875 | Rgy675);
assign L7a875 = (N8a875 & U8a875);
assign U8a875 = (Cg7875 | Kgy675);
assign N8a875 = (N29875 | Pfy675);
assign T4a875 = (~(H5a875 & Shm775));
assign Shm775 = (!Lwl775);
assign H5a875 = (Kw2875 & Rw2875);
assign Y3a875 = (~(hrdata_i[28] & Fy1875));
assign Fy8875 = (~(Aft775 & Sy1l85[12]));
assign Dx8875 = (Eg1875 & B9a875);
assign B9a875 = (~(vis_pc_o[11] & P60775));
assign Ygr675 = (~(I9a875 & P9a875));
assign P9a875 = (W9a875 & Daa875);
assign Daa875 = (~(E52l85[12] & Ykt775));
assign Ykt775 = (W60775 & O6v775);
assign W60775 = (F80775 & H90775);
assign W9a875 = (Kaa875 & Raa875);
assign Raa875 = (Vft775 | Bde775);
assign Bde775 = (Yaa875 & Fba875);
assign Fba875 = (Mba875 & Tba875);
assign Tba875 = (Pq0875 | Ve1875);
assign Ve1875 = (Nqz775 & Ua1875);
assign Ua1875 = (~(Aca875 & W41875));
assign Aca875 = (T5a775 & Kny675);
assign Nqz775 = (!Ijt775);
assign Ijt775 = (~(R67875 & Ga1875));
assign Ga1875 = (!Y67875);
assign Y67875 = (W41875 & C1g775);
assign R67875 = (Swl775 | W41875);
assign Pq0875 = (Hca875 & Oca875);
assign Oca875 = (Vca875 & Cda875);
assign Cda875 = (Ip1875 | Otm775);
assign Otm775 = (Jda875 & Qda875);
assign Qda875 = (Xda875 & Eea875);
assign Eea875 = (~(Eh7875 & Lea875));
assign Xda875 = (Jg7875 | Uey675);
assign Jda875 = (Sea875 & Zea875);
assign Zea875 = (Cg7875 | Ney675);
assign Sea875 = (Sh7875 | Gey675);
assign Vca875 = (~(Pp1875 & Gfa875));
assign Gfa875 = (~(Nfa875 & Ufa875));
assign Ufa875 = (Bga875 & Iga875);
assign Iga875 = (~(Pf2l85[5] & Wn4775));
assign Bga875 = (Pga875 & Wga875);
assign Wga875 = (~(st_calib_i[5] & Nv1875));
assign Pga875 = (~(V72l85[5] & Kn5775));
assign Nfa875 = (Dha875 & Kha875);
assign Kha875 = (~(Dx1875 & Gi2l85[5]));
assign Dha875 = (~(Iw1875 & Yg2l85[5]));
assign Hca875 = (Rha875 & Yha875);
assign Yha875 = (~(Yx1875 & Evm775));
assign Evm775 = (~(Fia875 & Mia875));
assign Mia875 = (Tia875 & Aja875);
assign Aja875 = (Jg7875 | Sdy675);
assign Tia875 = (Sh7875 | Nly675);
assign Fia875 = (Hja875 & Oja875);
assign Oja875 = (~(Eh7875 & Vja875));
assign Hja875 = (Cg7875 | Uly675);
assign Rha875 = (~(hrdata_i[5] & Fy1875));
assign Mba875 = (Rr0875 | Oe1875);
assign Oe1875 = (I41875 & Cka875);
assign Cka875 = (~(W41875 & Jka875));
assign Jka875 = (~(Qka875 & Xka875));
assign Xka875 = (~(Ela875 & O01875));
assign Ela875 = (~(Lla875 & Sla875));
assign Lla875 = (Zry675 | Vxo675);
assign Qka875 = (C4z675 & Za1775);
assign C4z675 = (Agl775 | Zry675);
assign Agl775 = (Xza775 | K1z675);
assign I41875 = (!Dlz775);
assign Dlz775 = (~(Zla875 & Nd5875));
assign Nd5875 = (~(W41875 & Gma875));
assign Gma875 = (~(Bvh675 & Nma875));
assign Nma875 = (~(Wxf775 & Uma875));
assign Uma875 = (Pw9775 | K1z675);
assign Zla875 = (Uwm775 | W41875);
assign Rr0875 = (Bna875 & Ina875);
assign Ina875 = (Pna875 & Wna875);
assign Wna875 = (Ip1875 | R6m775);
assign R6m775 = (Doa875 & Koa875);
assign Koa875 = (Roa875 & Yoa875);
assign Yoa875 = (~(Eh7875 & Fpa875));
assign Roa875 = (Sh7875 | Lky675);
assign Doa875 = (Mpa875 & Tpa875);
assign Tpa875 = (Cg7875 | Sky675);
assign Mpa875 = (Jg7875 | Zky675);
assign Pna875 = (~(Pp1875 & Aqa875));
assign Aqa875 = (~(Hqa875 & Oqa875));
assign Oqa875 = (Vqa875 & Cra875);
assign Cra875 = (~(V72l85[13] & Kn5775));
assign Vqa875 = (Jra875 & Qra875);
assign Qra875 = (~(Xqj775 & Ky1775));
assign Ky1775 = (~(Xra875 & Esa875));
assign Esa875 = (~(Lsa875 & Ssa875));
assign Lsa875 = (~(Zsa875 & I14875));
assign Zsa875 = (K42875 ? Nta875 : Gta875);
assign Nta875 = (Uta875 & Bua875);
assign Bua875 = (~(R42875 & Vk9875));
assign Uta875 = (F52875 ? Pua875 : Iua875);
assign Pua875 = (Wua875 | Dva875);
assign Iua875 = (Yva875 ? Rva875 : Kva875);
assign Gta875 = (Fwa875 & Mwa875);
assign Mwa875 = (Ql9875 ? Axa875 : Twa875);
assign Axa875 = (Hxa875 | Oxa875);
assign Twa875 = (Wo9875 | Vxa875);
assign Fwa875 = (Cya875 & Jya875);
assign Jya875 = (~(A62875 & Rp9875));
assign Cya875 = (~(T52875 & Bo9875));
assign Jra875 = (~(st_calib_i[13] & Nv1875));
assign Hqa875 = (Qya875 & Xya875);
assign Xya875 = (~(Iw1875 & Yg2l85[13]));
assign Qya875 = (Eza875 & Lza875);
assign Lza875 = (~(Pf2l85[13] & Wn4775));
assign Eza875 = (~(Dx1875 & Gi2l85[13]));
assign Bna875 = (Sza875 & Zza875);
assign Zza875 = (~(Yx1875 & J9m775));
assign J9m775 = (~(G0b875 & N0b875));
assign N0b875 = (U0b875 & B1b875);
assign B1b875 = (~(Eh7875 & I1b875));
assign U0b875 = (Sh7875 | Jjy675);
assign G0b875 = (P1b875 & W1b875);
assign W1b875 = (Cg7875 | Qjy675);
assign P1b875 = (Jg7875 | Xjy675);
assign Sza875 = (~(hrdata_i[13] & Fy1875));
assign Yaa875 = (D2b875 & K2b875);
assign K2b875 = (Bq0875 | Qf1875);
assign Qf1875 = (!Kj1875);
assign Kj1875 = (~(Z91875 & X81875));
assign X81875 = (~(W41875 & R2b875));
assign Z91875 = (~(Cb5875 & Ubm775));
assign Cb5875 = (Sc5875 & Z21875);
assign Bq0875 = (Y2b875 & F3b875);
assign F3b875 = (M3b875 & T3b875);
assign T3b875 = (Ip1875 | Ddm775);
assign Ddm775 = (A4b875 & H4b875);
assign H4b875 = (O4b875 & V4b875);
assign V4b875 = (~(Eh7875 & C5b875));
assign O4b875 = (Sh7875 | Aiy675);
assign A4b875 = (J5b875 & Q5b875);
assign Q5b875 = (Cg7875 | Hiy675);
assign J5b875 = (Jg7875 | Oiy675);
assign Ip1875 = (!Ob4875);
assign Ob4875 = (~(Nt3875 | Kll775));
assign M3b875 = (~(Pp1875 & X5b875));
assign X5b875 = (~(E6b875 & L6b875));
assign L6b875 = (S6b875 & Z6b875);
assign Z6b875 = (~(Pf2l85[21] & Wn4775));
assign S6b875 = (G7b875 & N7b875);
assign N7b875 = (~(st_calib_i[21] & Nv1875));
assign G7b875 = (~(V72l85[21] & Kn5775));
assign E6b875 = (U7b875 & B8b875);
assign B8b875 = (~(Dx1875 & Gi2l85[21]));
assign U7b875 = (~(Iw1875 & Yg2l85[21]));
assign Y2b875 = (I8b875 & P8b875);
assign P8b875 = (~(Yx1875 & Ofm775));
assign Ofm775 = (~(W8b875 & D9b875));
assign D9b875 = (K9b875 & R9b875);
assign R9b875 = (Jg7875 | Mhy675);
assign K9b875 = (~(Eh7875 & Y9b875));
assign W8b875 = (Fab875 & Mab875);
assign Mab875 = (Sh7875 | Ygy675);
assign Fab875 = (Cg7875 | Fhy675);
assign Yx1875 = (~(Nt3875 | Iqm775));
assign I8b875 = (~(hrdata_i[21] & Fy1875));
assign D2b875 = (Kr0875 | Xf1875);
assign Xf1875 = (!Yj1875);
assign Yj1875 = (~(Tab875 & Abb875));
assign Abb875 = (~(Hbb875 & Obb875));
assign Obb875 = (~(Zry675 | Vxo675));
assign Tab875 = (~(Tz0875 | Fz0875));
assign Fz0875 = (G31875 & Z21875);
assign Tz0875 = (Hbb875 & Vbb875);
assign Vbb875 = (~(Zh1775 | K1z675));
assign Hbb875 = (~(O01875 | Z21875));
assign Kr0875 = (Ccb875 & Jcb875);
assign Jcb875 = (Qcb875 & Xcb875);
assign Xcb875 = (~(Nl4875 & Gi2l85[29]));
assign Nl4875 = (Dx1875 & Pp1875);
assign Qcb875 = (Edb875 & Ek4875);
assign Ek4875 = (~(Ldb875 & Pp1875));
assign Ldb875 = (!N04875);
assign Edb875 = (~(hrdata_i[29] & Fy1875));
assign Ccb875 = (Sdb875 & Zdb875);
assign Zdb875 = (Lk4875 | Geb875);
assign Lk4875 = (~(Iw1875 & Pp1875));
assign Sdb875 = (~(Gu2875 & Neb875));
assign Neb875 = (~(Ueb875 & Bfb875));
assign Bfb875 = (Ifb875 | Lwl775);
assign Ueb875 = (~(Wqm775 & Pfb875));
assign Pfb875 = (Krm775 | Iqm775);
assign Krm775 = (~(Wfb875 & Dgb875));
assign Dgb875 = (Kgb875 & Rgb875);
assign Rgb875 = (Sh7875 | Ify675);
assign Kgb875 = (Jg7875 | Cjy675);
assign Wfb875 = (Ygb875 & Fhb875);
assign Fhb875 = (Cg7875 | Dgy675);
assign Ygb875 = (~(Eh7875 & Mhb875));
assign Wqm775 = (Thb875 & Ifb875);
assign Ifb875 = (~(Aib875 & Kw2875));
assign Aib875 = (Qj4875 ? Yw2875 : Rw2875);
assign Qj4875 = (Fx2875 & Sh7875);
assign Fx2875 = (~(Hib875 | Oib875));
assign Thb875 = (Hi4875 | Kll775);
assign Hi4875 = (~(Vib875 & Cjb875));
assign Cjb875 = (Jjb875 & Qjb875);
assign Qjb875 = (~(Eh7875 & Xjb875));
assign Jjb875 = (Sh7875 | Pfy675);
assign Vib875 = (Ekb875 & Lkb875);
assign Lkb875 = (Cg7875 | Wfy675);
assign Ekb875 = (Jg7875 | Kgy675);
assign Kaa875 = (~(Aft775 & Sy1l85[13]));
assign Aft775 = (~(P60775 | F80775));
assign I9a875 = (Eg1875 & Skb875);
assign Skb875 = (~(vis_pc_o[12] & P60775));
assign Eg1875 = (Oft775 & Zkb875);
assign Zkb875 = (Kse775 | Vft775);
assign Vft775 = (!Bi1875);
assign Bi1875 = (~(P60775 | H90775));
assign Kse775 = (~(C11875 & Glb875));
assign Glb875 = (~(Nlb875 & X11875));
assign X11875 = (~(Ulb875 & hresp_i));
assign Ulb875 = (Pp1875 & W41875);
assign Nlb875 = (!Bmb875);
assign Bmb875 = (W41875 ? Imb875 : Gim775);
assign W41875 = (!Z21875);
assign Z21875 = (~(Wbg775 & Pmb875));
assign Pmb875 = (~(Wmb875 & Af1775));
assign Wmb875 = (~(Wc1775 | X5p675));
assign Wbg775 = (!Dnb875);
assign Imb875 = (~(Knb875 & Rnb875));
assign Rnb875 = (~(Ynb875 & Zx6775));
assign Ynb875 = (~(Cm2775 | Mwo675));
assign Knb875 = (A2l775 | Xza775);
assign Gim775 = (!P5m775);
assign P5m775 = (B5m775 | G31875);
assign G31875 = (!Oul775);
assign Oul775 = (Rll775 | B41875);
assign Rll775 = (Fob875 | Mob875);
assign B5m775 = (~(N31875 & Swl775));
assign Swl775 = (~(Tob875 & Kkm775));
assign Kkm775 = (Fob875 & Apb875);
assign Fob875 = (!Hpb875);
assign Tob875 = (~(B41875 | Opb875));
assign N31875 = (Vpb875 & Uwm775);
assign Uwm775 = (~(Jvl775 & Ubm775));
assign Jvl775 = (Rkm775 & Flm775);
assign Vpb875 = (~(Sc5875 & Ubm775));
assign Ubm775 = (Y1z675 | Cqb875);
assign Sc5875 = (!Hul775);
assign Hul775 = (Onl775 | B41875);
assign B41875 = (!Flm775);
assign Flm775 = (~(Ezo675 & Jqb875));
assign Jqb875 = (~(Qhl775 & Xhl775));
assign Xhl775 = (Qqb875 | Xqb875);
assign Xqb875 = (X5y675 & Q5y675);
assign Qhl775 = (Erb875 & Lrb875);
assign Lrb875 = (~(Srb875 & Zrb875));
assign Zrb875 = (Gsb875 & Nsb875);
assign Nsb875 = (~(Xwi675 | Rto675));
assign Gsb875 = (~(Pui675 | Tvi675));
assign Srb875 = (Usb875 & Btb875);
assign Usb875 = (~(Hsi675 | Lti675));
assign Erb875 = (Qqb875 | E6y675);
assign Onl775 = (Apb875 | Hpb875);
assign Apb875 = (!Mob875);
assign C11875 = (~(Itb875 & Ptb875));
assign Ptb875 = (Wtb875 & Dub875);
assign Dub875 = (Kub875 | Epz775);
assign Epz775 = (Rub875 & Yub875);
assign Yub875 = (~(hrdata_i[15] & Fy1875));
assign Rub875 = (Fvb875 & Mvb875);
assign Mvb875 = (Nt3875 | Yll775);
assign Yll775 = (!Tvb875);
assign Tvb875 = (Kll775 ? Lhm775 : C9m775);
assign Lhm775 = (~(Awb875 & Hwb875));
assign Hwb875 = (Owb875 & Vwb875);
assign Vwb875 = (N29875 | Hiy675);
assign Owb875 = (Sh7875 | Oiy675);
assign Awb875 = (Cxb875 & Jxb875);
assign Jxb875 = (Cg7875 | Viy675);
assign Cxb875 = (Jg7875 | Jjy675);
assign C9m775 = (~(Qxb875 & Xxb875));
assign Xxb875 = (Eyb875 & Lyb875);
assign Lyb875 = (Cg7875 | Eky675);
assign Eky675 = (!Fpa875);
assign Fpa875 = (~(Syb875 & Zyb875));
assign Zyb875 = (Gzb875 & Nzb875);
assign Nzb875 = (Uzb875 & B0c875);
assign B0c875 = (~(I0c875 & vis_r0_o[16]));
assign Uzb875 = (~(P0c875 & vis_r2_o[16]));
assign Gzb875 = (W0c875 & D1c875);
assign D1c875 = (~(K1c875 & vis_r5_o[16]));
assign W0c875 = (~(R1c875 & vis_r4_o[16]));
assign Syb875 = (Y1c875 & F2c875);
assign F2c875 = (M2c875 & T2c875);
assign T2c875 = (~(A3c875 & vis_r7_o[16]));
assign M2c875 = (~(H3c875 & vis_r3_o[16]));
assign Y1c875 = (O3c875 & V3c875);
assign V3c875 = (~(C4c875 & vis_r1_o[16]));
assign O3c875 = (~(J4c875 & vis_r6_o[16]));
assign Eyb875 = (N29875 | Qjy675);
assign Qxb875 = (Q4c875 & X4c875);
assign X4c875 = (Sh7875 | Xjy675);
assign Q4c875 = (Jg7875 | Lky675);
assign Fvb875 = (~(Pp1875 & E5c875));
assign E5c875 = (~(L5c875 & S5c875));
assign S5c875 = (Z5c875 & G6c875);
assign G6c875 = (N6c875 & U6c875);
assign U6c875 = (B7c875 & S12875);
assign S12875 = (~(Opj775 & Bi8875));
assign B7c875 = (~(Rg5775 & Mb2l85[59]));
assign N6c875 = (I7c875 & P7c875);
assign P7c875 = (~(Fh5775 & Mb2l85[51]));
assign I7c875 = (~(Th5775 & Mb2l85[43]));
assign Z5c875 = (W7c875 & D8c875);
assign D8c875 = (K8c875 & R8c875);
assign R8c875 = (~(Hi5775 & Mb2l85[35]));
assign K8c875 = (~(Vi5775 & Mb2l85[27]));
assign W7c875 = (Y8c875 & F9c875);
assign F9c875 = (~(Jj5775 & Mb2l85[19]));
assign Y8c875 = (~(Xj5775 & Mb2l85[11]));
assign L5c875 = (M9c875 & T9c875);
assign T9c875 = (Aac875 & Hac875);
assign Hac875 = (Oac875 & Vac875);
assign Vac875 = (~(Lk5775 & Mb2l85[3]));
assign Oac875 = (~(S22775 & Xqj775));
assign S22775 = (B14875 & Cbc875);
assign Cbc875 = (~(Jbc875 & I14875));
assign Jbc875 = (Zd4875 ? Ql9875 : F52875);
assign B14875 = (!G22875);
assign G22875 = (~(Xra875 & Ssa875));
assign Xra875 = (~(Cep675 | Wcp675));
assign Aac875 = (Qbc875 & Xbc875);
assign Xbc875 = (~(st_calib_i[15] & Nv1875));
assign Qbc875 = (~(V72l85[15] & Kn5775));
assign M9c875 = (Ecc875 & Lcc875);
assign Lcc875 = (~(Iw1875 & Yg2l85[15]));
assign Ecc875 = (Scc875 & Zcc875);
assign Zcc875 = (~(Pf2l85[15] & Wn4775));
assign Scc875 = (~(Dx1875 & Gi2l85[15]));
assign Kub875 = (Gdc875 & Ndc875);
assign Ndc875 = (Jbk775 | Zry675);
assign Jbk775 = (D1z675 | Xza775);
assign Gdc875 = (~(Udc875 & O01875));
assign O01875 = (!M62l85[1]);
assign Wtb875 = (Bec875 & Lwl775);
assign Bec875 = (~(Iec875 & Qoz775));
assign Qoz775 = (~(Pec875 & Wec875));
assign Wec875 = (~(Pp1875 & Dfc875));
assign Dfc875 = (~(Kfc875 & Rfc875));
assign Rfc875 = (Yfc875 & Fgc875);
assign Fgc875 = (Mgc875 & Tgc875);
assign Tgc875 = (Ahc875 & Hhc875);
assign Hhc875 = (~(Rg5775 & Mb2l85[57]));
assign Ahc875 = (~(Fh5775 & Mb2l85[49]));
assign Mgc875 = (Ohc875 & Vhc875);
assign Vhc875 = (~(Th5775 & Mb2l85[41]));
assign Ohc875 = (~(Hi5775 & Mb2l85[33]));
assign Yfc875 = (Cic875 & Jic875);
assign Jic875 = (~(Xj5775 & Mb2l85[9]));
assign Cic875 = (Qic875 & Xic875);
assign Xic875 = (~(Vi5775 & Mb2l85[25]));
assign Qic875 = (~(Jj5775 & Mb2l85[17]));
assign Kfc875 = (Ejc875 & Ljc875);
assign Ljc875 = (Sjc875 & Zjc875);
assign Zjc875 = (~(V72l85[7] & Kn5775));
assign Sjc875 = (Gkc875 & Nkc875);
assign Nkc875 = (~(Lk5775 & Mb2l85[1]));
assign Gkc875 = (~(st_calib_i[7] & Nv1875));
assign Ejc875 = (Ukc875 & Blc875);
assign Blc875 = (~(Iw1875 & Yg2l85[7]));
assign Ukc875 = (Ilc875 & Plc875);
assign Plc875 = (~(Pf2l85[7] & Wn4775));
assign Ilc875 = (~(Dx1875 & Gi2l85[7]));
assign Pec875 = (Wlc875 & Dmc875);
assign Dmc875 = (Nt3875 | Hnl775);
assign Hnl775 = (Iqm775 ? Xum775 : Lam775);
assign Xum775 = (Kmc875 & Rmc875);
assign Rmc875 = (Ymc875 & Fnc875);
assign Fnc875 = (Sh7875 | Sdy675);
assign Sdy675 = (!Jn7875);
assign Jn7875 = (~(Mnc875 & Tnc875));
assign Tnc875 = (Aoc875 & Hoc875);
assign Hoc875 = (Ooc875 & Voc875);
assign Voc875 = (~(I0c875 & vis_r0_o[9]));
assign Ooc875 = (~(P0c875 & vis_r2_o[9]));
assign Aoc875 = (Cpc875 & Jpc875);
assign Jpc875 = (~(K1c875 & vis_r5_o[9]));
assign Cpc875 = (~(R1c875 & vis_r4_o[9]));
assign Mnc875 = (Qpc875 & Xpc875);
assign Xpc875 = (Eqc875 & Lqc875);
assign Lqc875 = (~(A3c875 & vis_r7_o[9]));
assign Eqc875 = (~(H3c875 & vis_r3_o[9]));
assign Qpc875 = (Sqc875 & Zqc875);
assign Zqc875 = (~(C4c875 & vis_r1_o[9]));
assign Sqc875 = (~(J4c875 & vis_r6_o[9]));
assign Ymc875 = (Cg7875 | Zdy675);
assign Zdy675 = (!Lea875);
assign Lea875 = (~(Grc875 & Nrc875));
assign Nrc875 = (Urc875 & Bsc875);
assign Bsc875 = (Isc875 & Psc875);
assign Psc875 = (~(I0c875 & vis_r0_o[8]));
assign Isc875 = (~(P0c875 & vis_r2_o[8]));
assign Urc875 = (Wsc875 & Dtc875);
assign Dtc875 = (~(K1c875 & vis_r5_o[8]));
assign Wsc875 = (~(R1c875 & vis_r4_o[8]));
assign Grc875 = (Ktc875 & Rtc875);
assign Rtc875 = (Ytc875 & Fuc875);
assign Fuc875 = (~(A3c875 & vis_r7_o[8]));
assign Ytc875 = (~(H3c875 & vis_r3_o[8]));
assign Ktc875 = (Muc875 & Tuc875);
assign Tuc875 = (~(C4c875 & vis_r1_o[8]));
assign Muc875 = (~(J4c875 & vis_r6_o[8]));
assign Kmc875 = (Avc875 & Hvc875);
assign Hvc875 = (N29875 | Uly675);
assign Avc875 = (Jg7875 | Gey675);
assign Lam775 = (Ovc875 & Vvc875);
assign Vvc875 = (Cwc875 & Jwc875);
assign Jwc875 = (Jg7875 | Nly675);
assign Nly675 = (Qwc875 & Xwc875);
assign Xwc875 = (Exc875 & Lxc875);
assign Lxc875 = (Sxc875 & Zxc875);
assign Zxc875 = (~(I0c875 & vis_r0_o[11]));
assign Sxc875 = (~(P0c875 & vis_r2_o[11]));
assign Exc875 = (Gyc875 & Nyc875);
assign Nyc875 = (~(K1c875 & vis_r5_o[11]));
assign Gyc875 = (~(R1c875 & vis_r4_o[11]));
assign Qwc875 = (Uyc875 & Bzc875);
assign Bzc875 = (Izc875 & Pzc875);
assign Pzc875 = (~(A3c875 & vis_r7_o[11]));
assign Izc875 = (~(H3c875 & vis_r3_o[11]));
assign Uyc875 = (Wzc875 & D0d875);
assign D0d875 = (~(C4c875 & vis_r1_o[11]));
assign Wzc875 = (~(J4c875 & vis_r6_o[11]));
assign Cwc875 = (Cg7875 | Gly675);
assign Gly675 = (!Vja875);
assign Vja875 = (~(K0d875 & R0d875));
assign R0d875 = (Y0d875 & F1d875);
assign F1d875 = (M1d875 & T1d875);
assign T1d875 = (~(I0c875 & vis_r0_o[12]));
assign M1d875 = (~(P0c875 & vis_r2_o[12]));
assign Y0d875 = (A2d875 & H2d875);
assign H2d875 = (~(K1c875 & vis_r5_o[12]));
assign A2d875 = (~(R1c875 & vis_r4_o[12]));
assign K0d875 = (O2d875 & V2d875);
assign V2d875 = (C3d875 & J3d875);
assign J3d875 = (~(A3c875 & vis_r7_o[12]));
assign C3d875 = (~(H3c875 & vis_r3_o[12]));
assign O2d875 = (Q3d875 & X3d875);
assign X3d875 = (~(C4c875 & vis_r1_o[12]));
assign Q3d875 = (~(J4c875 & vis_r6_o[12]));
assign Ovc875 = (E4d875 & L4d875);
assign L4d875 = (N29875 | Sky675);
assign E4d875 = (Sh7875 | Zky675);
assign Wlc875 = (~(hrdata_i[7] & Fy1875));
assign Iec875 = (~(A2l775 & S4d875));
assign S4d875 = (~(Z4d875 & Xza775));
assign Z4d875 = (~(K1z675 & G5d875));
assign G5d875 = (M62l85[0] | M62l85[1]);
assign A2l775 = (!Ytr775);
assign Itb875 = (N5d875 & U5d875);
assign U5d875 = (~(M62l85[1] & B6d875));
assign B6d875 = (~(I6d875 & P6d875));
assign P6d875 = (~(W6d875 & V0g775));
assign W6d875 = (~(Gqz775 | M62l85[0]));
assign Gqz775 = (D7d875 & K7d875);
assign K7d875 = (~(Pp1875 & R7d875));
assign R7d875 = (~(Y7d875 & F8d875));
assign F8d875 = (M8d875 & T8d875);
assign T8d875 = (A9d875 & H9d875);
assign H9d875 = (O9d875 & V9d875);
assign V9d875 = (~(Bm5775 & C92l85[1]));
assign O9d875 = (~(Rg5775 & Mb2l85[61]));
assign A9d875 = (Cad875 & Jad875);
assign Jad875 = (~(Fh5775 & Mb2l85[53]));
assign Cad875 = (~(Th5775 & Mb2l85[45]));
assign M8d875 = (Qad875 & Xad875);
assign Xad875 = (~(Jj5775 & Mb2l85[21]));
assign Qad875 = (Ebd875 & Lbd875);
assign Lbd875 = (~(Hi5775 & Mb2l85[37]));
assign Ebd875 = (~(Vi5775 & Mb2l85[29]));
assign Y7d875 = (Sbd875 & Zbd875);
assign Zbd875 = (Gcd875 & Ncd875);
assign Ncd875 = (Ucd875 & Bdd875);
assign Bdd875 = (~(Xj5775 & Mb2l85[13]));
assign Ucd875 = (~(Lk5775 & Mb2l85[5]));
assign Gcd875 = (Idd875 & Pdd875);
assign Pdd875 = (~(st_calib_i[23] & Nv1875));
assign Idd875 = (~(V72l85[23] & Kn5775));
assign Kn5775 = (~(Wdd875 | Ded875));
assign Sbd875 = (Ked875 & Red875);
assign Red875 = (~(Iw1875 & Yg2l85[23]));
assign Ked875 = (Yed875 & Ffd875);
assign Ffd875 = (~(Pf2l85[23] & Wn4775));
assign Wn4775 = (~(Wj7875 | Ii8875));
assign Yed875 = (~(Dx1875 & Gi2l85[23]));
assign D7d875 = (Mfd875 & Tfd875);
assign Tfd875 = (Nt3875 | Anl775);
assign Anl775 = (Kll775 ? Bw8875 : Vfm775);
assign Bw8875 = (Agd875 & Hgd875);
assign Hgd875 = (Ogd875 & Vgd875);
assign Vgd875 = (N29875 | Wfy675);
assign Ogd875 = (Sh7875 | Kgy675);
assign Agd875 = (Chd875 & Jhd875);
assign Jhd875 = (~(Hib875 & Qhd875));
assign Chd875 = (~(Oib875 & Y9b875));
assign Vfm775 = (Xhd875 & Eid875);
assign Eid875 = (Lid875 & Sid875);
assign Sid875 = (Sh7875 | Mhy675);
assign Mhy675 = (!U38875);
assign U38875 = (~(Zid875 & Gjd875));
assign Gjd875 = (Njd875 & Ujd875);
assign Ujd875 = (Bkd875 & Ikd875);
assign Ikd875 = (~(I0c875 & vis_r0_o[25]));
assign Bkd875 = (~(P0c875 & vis_r2_o[25]));
assign Njd875 = (Pkd875 & Wkd875);
assign Wkd875 = (~(K1c875 & vis_r5_o[25]));
assign Pkd875 = (~(R1c875 & vis_r4_o[25]));
assign Zid875 = (Dld875 & Kld875);
assign Kld875 = (Rld875 & Yld875);
assign Yld875 = (~(A3c875 & vis_r7_o[25]));
assign Rld875 = (~(H3c875 & vis_r3_o[25]));
assign Dld875 = (Fmd875 & Mmd875);
assign Mmd875 = (~(C4c875 & vis_r1_o[25]));
assign Fmd875 = (~(J4c875 & vis_r6_o[25]));
assign Lid875 = (N29875 | Fhy675);
assign Xhd875 = (Tmd875 & And875);
assign And875 = (Cg7875 | Thy675);
assign Tmd875 = (Jg7875 | Aiy675);
assign Mfd875 = (~(hrdata_i[23] & Fy1875));
assign I6d875 = (~(Udc875 & Zpz775));
assign Zpz775 = (~(Hnd875 & Ond875));
assign Ond875 = (~(Pp1875 & Vnd875));
assign Vnd875 = (~(Cod875 & Jod875));
assign Jod875 = (Qod875 & Xod875);
assign Xod875 = (Epd875 & Lpd875);
assign Lpd875 = (Spd875 & N04875);
assign Spd875 = (~(Nl5775 & Ha2l85[1]));
assign Nl5775 = (Zpd875 & Ar3775);
assign Epd875 = (Gqd875 & Nqd875);
assign Nqd875 = (~(Bm5775 & Ge2l85[1]));
assign Bm5775 = (Uqd875 & Brd875);
assign Uqd875 = (~(F59875 | Ilz675));
assign Gqd875 = (~(Rg5775 & Mb2l85[63]));
assign Rg5775 = (~(Ird875 | Wj7875));
assign Qod875 = (Prd875 & Wrd875);
assign Wrd875 = (Dsd875 & Ksd875);
assign Ksd875 = (~(Fh5775 & Mb2l85[55]));
assign Fh5775 = (~(Ded875 | Wj7875));
assign Wj7875 = (~(Toj775 & Ilz675));
assign Dsd875 = (~(Th5775 & Mb2l85[47]));
assign Th5775 = (~(Wdd875 | Ii8875));
assign Prd875 = (Rsd875 & Ysd875);
assign Ysd875 = (~(Hi5775 & Mb2l85[39]));
assign Hi5775 = (~(Wdd875 | Hr3775));
assign Hr3775 = (!Y49875);
assign Rsd875 = (~(Vi5775 & Mb2l85[31]));
assign Vi5775 = (Ftd875 & Zpd875);
assign Cod875 = (Mtd875 & Ttd875);
assign Ttd875 = (Aud875 & Hud875);
assign Hud875 = (Oud875 & Vud875);
assign Vud875 = (~(Jj5775 & Mb2l85[23]));
assign Jj5775 = (Ftd875 & Brd875);
assign Brd875 = (!Ded875);
assign Ded875 = (~(Ycr675 & Hhz675));
assign Ftd875 = (Toj775 & Aar675);
assign Oud875 = (~(Xj5775 & Mb2l85[15]));
assign Xj5775 = (~(Cvd875 | Apj775));
assign Aud875 = (Jvd875 & Qvd875);
assign Qvd875 = (~(Lk5775 & Mb2l85[7]));
assign Lk5775 = (~(Cvd875 | Bn4775));
assign Jvd875 = (~(Wcp675 & Xqj775));
assign Xqj775 = (~(Apj775 | F59875));
assign F59875 = (!Bi8875);
assign Bi8875 = (~(Sjz675 | O8r675));
assign Mtd875 = (Xvd875 & Ewd875);
assign Ewd875 = (~(Iw1875 & Yg2l85[31]));
assign Iw1875 = (Nm4775 & Lwd875);
assign Xvd875 = (Swd875 & Zwd875);
assign Zwd875 = (~(st_calib_i[25] & Nv1875));
assign Nv1875 = (~(Wdd875 | Ird875));
assign Wdd875 = (Cvd875 | Aar675);
assign Cvd875 = (G6z675 | Sjz675);
assign Sjz675 = (!Mbr675);
assign Swd875 = (~(Dx1875 & Gi2l85[31]));
assign Dx1875 = (Toj775 & Lwd875);
assign Lwd875 = (~(Apj775 & Bn4775));
assign Bn4775 = (!Opj775);
assign Opj775 = (Y49875 & Aar675);
assign Apj775 = (Ilz675 | Ii8875);
assign Ii8875 = (Hhz675 | Ycr675);
assign Hhz675 = (!Ker675);
assign Toj775 = (~(G6z675 | Mbr675));
assign G6z675 = (!O8r675);
assign Hnd875 = (Gxd875 & Nxd875);
assign Nxd875 = (Nt3875 | Cvl775);
assign Cvl775 = (Byd875 ? Lwl775 : Uxd875);
assign Byd875 = (Iyd875 & Kw2875);
assign Kw2875 = (Ezo675 & Jj4875);
assign Jj4875 = (~(Cj4875 & Kll775));
assign Iyd875 = (Jg7875 ? Yw2875 : Rw2875);
assign Rw2875 = (~(Iqm775 & Yw2875));
assign Yw2875 = (!Cj4875);
assign Cj4875 = (Pyd875 & Mtl775);
assign Mtl775 = (!Opb875);
assign Opb875 = (K7s775 & Y1z675);
assign Pyd875 = (!Cqb875);
assign Cqb875 = (Wyd875 & Hib875);
assign Wyd875 = (~(Kll775 | Pkl775));
assign Pkl775 = (!Rkm775);
assign Rkm775 = (Mob875 & Hpb875);
assign Hpb875 = (Rto675 ? Kzd875 : Dzd875);
assign Kzd875 = (~(Rzd875 & Yzd875));
assign Rzd875 = (~(F0e875 & M0e875));
assign Dzd875 = (!F0e875);
assign Mob875 = (Rto675 ? A1e875 : T0e875);
assign A1e875 = (H1e875 | Jhl775);
assign Jhl775 = (~(Yzd875 | O1e875));
assign H1e875 = (O1e875 & Yzd875);
assign Yzd875 = (M0e875 | F0e875);
assign F0e875 = (~(V1e875 & C2e875));
assign C2e875 = (Qqb875 | S6y675);
assign V1e875 = (~(Btb875 & Tvi675));
assign O1e875 = (!T0e875);
assign T0e875 = (J2e875 & Q2e875);
assign Q2e875 = (Qqb875 | L6y675);
assign J2e875 = (~(Btb875 & Xwi675));
assign Kll775 = (!Iqm775);
assign Lwl775 = (~(X2e875 & C4i675));
assign X2e875 = (~(Wrl775 | Pfy675));
assign Wrl775 = (Rxg775 & E3e875);
assign E3e875 = (Bbg775 | Rto675);
assign Uxd875 = (Iqm775 ? Wkl775 : Dll775);
assign Iqm775 = (Rto675 ? S3e875 : L3e875);
assign S3e875 = (~(Z3e875 & M0e875));
assign M0e875 = (G4e875 | N4e875);
assign Z3e875 = (~(N4e875 & G4e875));
assign L3e875 = (!G4e875);
assign G4e875 = (~(U4e875 & B5e875));
assign B5e875 = (Qqb875 | N7y675);
assign U4e875 = (~(Btb875 & Pui675));
assign Wkl775 = (I5e875 & P5e875);
assign P5e875 = (W5e875 & D6e875);
assign D6e875 = (N29875 | Dgy675);
assign Dgy675 = (K6e875 & R6e875);
assign R6e875 = (Y6e875 & F7e875);
assign F7e875 = (M7e875 & T7e875);
assign T7e875 = (~(I0c875 & vis_r0_o[2]));
assign M7e875 = (~(P0c875 & vis_r2_o[2]));
assign Y6e875 = (A8e875 & H8e875);
assign H8e875 = (~(K1c875 & vis_r5_o[2]));
assign A8e875 = (~(R1c875 & vis_r4_o[2]));
assign K6e875 = (O8e875 & V8e875);
assign V8e875 = (C9e875 & J9e875);
assign J9e875 = (~(A3c875 & vis_r7_o[2]));
assign C9e875 = (~(H3c875 & vis_r3_o[2]));
assign O8e875 = (Q9e875 & X9e875);
assign X9e875 = (~(C4c875 & vis_r1_o[2]));
assign Q9e875 = (~(J4c875 & vis_r6_o[2]));
assign W5e875 = (Cg7875 | Bmy675);
assign I5e875 = (Eae875 & Lae875);
assign Lae875 = (Jg7875 | Pfy675);
assign Eae875 = (Sh7875 | Cjy675);
assign Dll775 = (Sae875 & Zae875);
assign Zae875 = (Gbe875 & Nbe875);
assign Nbe875 = (N29875 | Ney675);
assign N29875 = (!Eh7875);
assign Eh7875 = (~(Ube875 | Bce875));
assign Gbe875 = (Cg7875 | Bfy675);
assign Cg7875 = (!Oib875);
assign Oib875 = (Ube875 & Ice875);
assign Sae875 = (Pce875 & Wce875);
assign Wce875 = (Jg7875 | Ify675);
assign Ify675 = (!Q6a875);
assign Q6a875 = (~(Dde875 & Kde875));
assign Kde875 = (Rde875 & Yde875);
assign Yde875 = (Fee875 & Mee875);
assign Mee875 = (~(I0c875 & vis_r0_o[3]));
assign Fee875 = (~(P0c875 & vis_r2_o[3]));
assign Rde875 = (Tee875 & Afe875);
assign Afe875 = (~(K1c875 & vis_r5_o[3]));
assign Tee875 = (~(R1c875 & vis_r4_o[3]));
assign Dde875 = (Hfe875 & Ofe875);
assign Ofe875 = (Vfe875 & Cge875);
assign Cge875 = (~(A3c875 & vis_r7_o[3]));
assign Vfe875 = (~(H3c875 & vis_r3_o[3]));
assign Hfe875 = (Jge875 & Qge875);
assign Qge875 = (~(C4c875 & vis_r1_o[3]));
assign Jge875 = (~(J4c875 & vis_r6_o[3]));
assign Jg7875 = (!Hib875);
assign Hib875 = (Ube875 & Bce875);
assign Pce875 = (Sh7875 | Uey675);
assign Sh7875 = (Ice875 | Ube875);
assign Ube875 = (Rto675 ? Ehe875 : Xge875);
assign Ehe875 = (~(Lhe875 & N4e875));
assign N4e875 = (~(Xge875 & Bce875));
assign Lhe875 = (Bce875 | Xge875);
assign Bce875 = (!Ice875);
assign Xge875 = (She875 & Zhe875);
assign Zhe875 = (Qqb875 | May675);
assign She875 = (~(Btb875 & Lti675));
assign Ice875 = (~(Gie875 & Nie875));
assign Nie875 = (Qqb875 | Ldy675);
assign Qqb875 = (Nsj775 | Veg775);
assign Gie875 = (~(Btb875 & Hsi675));
assign Btb875 = (~(Nsj775 | L2g775));
assign Nsj775 = (!C4i675);
assign Nt3875 = (!Gu2875);
assign Gu2875 = (C4i675 & Uie875);
assign Uie875 = (~(Bje875 & Ije875));
assign Ije875 = (K1z675 | Zck775);
assign Bje875 = (~(Dnb875 | Ytr775));
assign Dnb875 = (D1z675 & Cg8775);
assign Gxd875 = (~(hrdata_i[31] & Fy1875));
assign Fy1875 = (Pje875 & Ar3775);
assign Ar3775 = (Nm4775 & Ilz675);
assign Ilz675 = (!Aar675);
assign Pje875 = (Pp1875 & Y49875);
assign Y49875 = (~(Ycr675 | Ker675));
assign Udc875 = (~(Wje875 & Sla875));
assign Sla875 = (Ryf775 | Mwo675);
assign Wje875 = (~(M62l85[0] & V0g775));
assign N5d875 = (~(hresp_i & Pp1875));
assign Pp1875 = (C4i675 & Dke875);
assign Dke875 = (~(Kke875 & Rke875));
assign Rke875 = (Vxo675 ? Zh1775 : Yke875);
assign Zh1775 = (!Waa775);
assign Waa775 = (Zck775 & Q91775);
assign Yke875 = (Af1775 | D1z675);
assign Af1775 = (!Gwf775);
assign Kke875 = (Fle875 & Cg8775);
assign Fle875 = (Yaw775 | Bvh675);
assign Oft775 = (~(O6v775 & Mle875));
assign Mle875 = (~(Tle875 & Ame875));
assign Ame875 = (~(Tth675 & Erj775));
assign Tle875 = (Hme875 & L40775);
assign Hme875 = (~(Lsh675 & C37775));
assign O6v775 = (!P60775);
assign P60775 = (Lcz675 | Fg5875);
assign Rgr675 = (~(Ome875 & Vme875));
assign Vme875 = (~(Zmo675 & Cne875));
assign Cne875 = (Prz775 | Lcz675);
assign Ome875 = (Jne875 | Lcz675);
assign Kgr675 = (Lcz675 ? Uhp675 : Qne875);
assign Lcz675 = (!hready_i);
assign Qne875 = (Xne875 & Eoe875);
assign Eoe875 = (Loe875 & Soe875);
assign Soe875 = (~(Zoe875 & Hph675));
assign Zoe875 = (~(Bwg775 | Rxg775));
assign Rxg775 = (!Gvg775);
assign Loe875 = (~(Gpe875 & Jqh675));
assign Gpe875 = (W1p675 & Npe875);
assign Npe875 = (~(Upe875 & Bqe875));
assign Upe875 = (~(Pw9775 & Iqe875));
assign Iqe875 = (V7g775 | Kxg775);
assign Kxg775 = (!Mch775);
assign V7g775 = (X5p675 & Mwo675);
assign Xne875 = (Qbz675 & Pqe875);
assign Pqe875 = (~(Svt775 & Wqe875));
assign Wqe875 = (Bqe875 | U50775);
assign Svt775 = (~(R2b875 & Uvg775));
assign Uvg775 = (~(Dre875 & Kre875));
assign Kre875 = (~(Rre875 & Yre875));
assign Yre875 = (~(Bvh675 | O4p675));
assign Rre875 = (~(Ycu775 | Lrh675));
assign Dre875 = (~(Fse875 & Cut775));
assign Qbz675 = (!Ts1775);
assign Ts1775 = (~(Abx775 & Mse875));
assign Mse875 = (~(Tse875 & Obx775));
assign Obx775 = (Ssa875 & Ate875);
assign Ate875 = (~(Hte875 & Ote875));
assign Ote875 = (Vte875 | Cue875);
assign Vte875 = (Xue875 ? Que875 : Jue875);
assign Hte875 = (Eve875 & Lve875);
assign Eve875 = (~(Sve875 & Zve875));
assign Zve875 = (B32875 ? Nwe875 : Gwe875);
assign Nwe875 = (~(Uwe875 | Bxe875));
assign Bxe875 = (~(Ixe875 | Pxe875));
assign Gwe875 = (~(Cue875 & Que875));
assign Sve875 = (Wxe875 & Dye875);
assign Wxe875 = (~(Kye875 & Xue875));
assign Ssa875 = (~(I14875 & Rye875));
assign I14875 = (P32875 & Xue875);
assign Xue875 = (!B32875);
assign B32875 = (Yye875 & Fze875);
assign Fze875 = (~(Mze875 & Tze875));
assign Tze875 = (~(A0f875 & H0f875));
assign H0f875 = (~(O0f875 & Uwe875));
assign Uwe875 = (U22875 ? Ha2l85[0] : C92l85[0]);
assign O0f875 = (~(Kye875 | V0f875));
assign V0f875 = (Ixe875 & Que875);
assign Kye875 = (P32875 ? C1f875 : Ge2l85[0]);
assign A0f875 = (Que875 | Ixe875);
assign Ixe875 = (!Jue875);
assign Jue875 = (U22875 ? Ha2l85[1] : C92l85[1]);
assign Que875 = (P32875 ? J1f875 : Ge2l85[1]);
assign Mze875 = (~(Rye875 & P32875));
assign Rye875 = (!Xe9875);
assign Yye875 = (Ifp675 | U22875);
assign U22875 = (Ogp675 & Q1f875);
assign Q1f875 = (~(X1f875 & Ifp675));
assign X1f875 = (E2f875 & L2f875);
assign L2f875 = (~(S2f875 & Z2f875));
assign Z2f875 = (G3f875 | C92l85[1]);
assign S2f875 = (N3f875 | C92l85[0]);
assign E2f875 = (~(C92l85[1] & G3f875));
assign P32875 = (~(E7r675 & U3f875));
assign U3f875 = (~(B4f875 & I4f875));
assign I4f875 = (~(J1f875 & Ycgk85));
assign B4f875 = (Xe9875 & Fdgk85);
assign Fdgk85 = (~(Mdgk85 & Tdgk85));
assign Tdgk85 = (~(Aegk85 & Ge2l85[0]));
assign Aegk85 = (!C1f875);
assign C1f875 = (K42875 ? Oegk85 : Hegk85);
assign Mdgk85 = (J1f875 | Ycgk85);
assign Ycgk85 = (!Ge2l85[1]);
assign J1f875 = (K42875 ? Cfgk85 : Vegk85);
assign K42875 = (!Zd4875);
assign Xe9875 = (~(Jfgk85 & A62875));
assign Jfgk85 = (Qfgk85 & Zd4875);
assign Zd4875 = (~(Xfgk85 & Eggk85));
assign Eggk85 = (Lggk85 | Sggk85);
assign Lggk85 = (F52875 | M52875);
assign Xfgk85 = (~(Zggk85 & Ghgk85));
assign Ghgk85 = (~(Vegk85 & Nhgk85));
assign Zggk85 = (Uhgk85 & Bigk85);
assign Bigk85 = (~(Iigk85 & Pigk85));
assign Pigk85 = (Nhgk85 | Vegk85);
assign Vegk85 = (Kjgk85 ? Djgk85 : Wigk85);
assign Nhgk85 = (!Cfgk85);
assign Cfgk85 = (F52875 ? Yjgk85 : Rjgk85);
assign Iigk85 = (Hegk85 | Fkgk85);
assign Fkgk85 = (!Oegk85);
assign Oegk85 = (~(Mkgk85 & Tkgk85));
assign Tkgk85 = (~(R42875 & Algk85));
assign Algk85 = (~(Hlgk85 & Olgk85));
assign R42875 = (F52875 & Wua875);
assign Mkgk85 = (F52875 ? Cmgk85 : Vlgk85);
assign F52875 = (!Gg9875);
assign Gg9875 = (~(Jmgk85 & Qmgk85));
assign Qmgk85 = (~(Xmgk85 & Engk85));
assign Engk85 = (~(Lngk85 & Sngk85));
assign Sngk85 = (~(Zngk85 & Gogk85));
assign Gogk85 = (Nogk85 & Uogk85);
assign Nogk85 = (~(Rjgk85 & Bpgk85));
assign Zngk85 = (~(Ipgk85 | Ppgk85));
assign Ppgk85 = (M52875 & Wpgk85);
assign Ipgk85 = (Fj9875 ? Kqgk85 : Dqgk85);
assign Lngk85 = (Bpgk85 | Rjgk85);
assign Rjgk85 = (M52875 ? Yqgk85 : Rqgk85);
assign Bpgk85 = (!Yjgk85);
assign Yjgk85 = (Fj9875 ? Mrgk85 : Frgk85);
assign Xmgk85 = (Sggk85 | M52875);
assign Jmgk85 = (~(Trgk85 & Asgk85));
assign Asgk85 = (~(Fj9875 | Hsgk85));
assign Fj9875 = (!Wua875);
assign Trgk85 = (~(Osgk85 | Vsgk85));
assign Cmgk85 = (Wua875 | Kqgk85);
assign Wua875 = (~(Ctgk85 & Jtgk85));
assign Jtgk85 = (~(Qtgk85 & Xtgk85));
assign Qtgk85 = (~(Eugk85 | Dva875));
assign Ctgk85 = (~(Lugk85 & Sugk85));
assign Sugk85 = (~(Zugk85 & Ok9875));
assign Ok9875 = (!Osgk85);
assign Zugk85 = (~(Vsgk85 | Hsgk85));
assign Lugk85 = (~(Gvgk85 & Nvgk85));
assign Nvgk85 = (~(Uvgk85 & Dqgk85));
assign Dqgk85 = (Hlgk85 & Olgk85);
assign Olgk85 = (~(Hsgk85 & Bwgk85));
assign Hlgk85 = (~(Iwgk85 & Vk9875));
assign Uvgk85 = (~(Kqgk85 | Pwgk85));
assign Pwgk85 = (~(Wwgk85 | Mrgk85));
assign Kqgk85 = (Dva875 ? Kxgk85 : Dxgk85);
assign Kxgk85 = (!Rxgk85);
assign Gvgk85 = (~(Mrgk85 & Wwgk85));
assign Wwgk85 = (!Frgk85);
assign Frgk85 = (Hsgk85 ? Fygk85 : Yxgk85);
assign Hsgk85 = (!Vk9875);
assign Vk9875 = (~(Mygk85 & Tygk85));
assign Tygk85 = (~(Azgk85 & Hzgk85));
assign Hzgk85 = (~(Ozgk85 & Vzgk85));
assign Vzgk85 = (~(C0hk85 & Bwgk85));
assign Bwgk85 = (Hk9875 ? Mb2l85[10] : Mb2l85[8]);
assign C0hk85 = (~(Iwgk85 | J0hk85));
assign J0hk85 = (Yxgk85 & Q0hk85);
assign Iwgk85 = (Osgk85 ? Mb2l85[12] : Mb2l85[14]);
assign Ozgk85 = (Q0hk85 | Yxgk85);
assign Q0hk85 = (!Fygk85);
assign Azgk85 = (Osgk85 | Vsgk85);
assign Mygk85 = (~(Hk9875 & X0hk85));
assign X0hk85 = (~(Yg2l85[5] & Gi2l85[5]));
assign Fygk85 = (Hk9875 ? Mb2l85[11] : Mb2l85[9]);
assign Hk9875 = (~(E1hk85 & Yg2l85[4]));
assign E1hk85 = (Gi2l85[4] & L1hk85);
assign L1hk85 = (~(S1hk85 & Yg2l85[5]));
assign S1hk85 = (Gi2l85[5] & Z1hk85);
assign Z1hk85 = (~(G2hk85 & N2hk85));
assign N2hk85 = (~(U2hk85 & Mb2l85[8]));
assign U2hk85 = (~(B3hk85 | Mb2l85[10]));
assign B3hk85 = (~(I3hk85 | Mb2l85[9]));
assign G2hk85 = (~(Mb2l85[9] & I3hk85));
assign Yxgk85 = (Osgk85 ? Mb2l85[13] : Mb2l85[15]);
assign Osgk85 = (P3hk85 & Yg2l85[6]);
assign P3hk85 = (Gi2l85[6] & W3hk85);
assign W3hk85 = (~(Vsgk85 & D4hk85));
assign D4hk85 = (~(K4hk85 & R4hk85));
assign R4hk85 = (~(Y4hk85 & Mb2l85[12]));
assign Y4hk85 = (~(F5hk85 | Mb2l85[14]));
assign F5hk85 = (~(M5hk85 | Mb2l85[13]));
assign K4hk85 = (~(Mb2l85[13] & M5hk85));
assign Vsgk85 = (Yg2l85[7] & Gi2l85[7]);
assign Mrgk85 = (Dva875 ? A6hk85 : T5hk85);
assign Dva875 = (!Ak9875);
assign Ak9875 = (~(H6hk85 & O6hk85));
assign O6hk85 = (~(V6hk85 & C7hk85));
assign C7hk85 = (~(J7hk85 & Q7hk85));
assign Q7hk85 = (~(X7hk85 & Rxgk85));
assign Rxgk85 = (Mj9875 ? Mb2l85[2] : Mb2l85[0]);
assign X7hk85 = (Dxgk85 & E8hk85);
assign E8hk85 = (L8hk85 | A6hk85);
assign Dxgk85 = (Tj9875 ? Z8hk85 : S8hk85);
assign J7hk85 = (~(A6hk85 & L8hk85));
assign V6hk85 = (~(Xtgk85 & Tj9875));
assign Tj9875 = (!Eugk85);
assign Xtgk85 = (~(Yg2l85[3] & Gi2l85[3]));
assign H6hk85 = (~(Mj9875 & G9hk85));
assign G9hk85 = (~(Yg2l85[1] & Gi2l85[1]));
assign A6hk85 = (Mj9875 ? Mb2l85[3] : Mb2l85[1]);
assign Mj9875 = (~(N9hk85 & Yg2l85[0]));
assign N9hk85 = (Gi2l85[0] & U9hk85);
assign U9hk85 = (~(Bahk85 & Yg2l85[1]));
assign Bahk85 = (Gi2l85[1] & Iahk85);
assign Iahk85 = (~(Pahk85 & Wahk85));
assign Wahk85 = (~(Dbhk85 & Mb2l85[0]));
assign Dbhk85 = (~(Kbhk85 | Mb2l85[2]));
assign Kbhk85 = (~(Rbhk85 | Mb2l85[1]));
assign Pahk85 = (~(Mb2l85[1] & Rbhk85));
assign T5hk85 = (!L8hk85);
assign L8hk85 = (Eugk85 ? Fchk85 : Ybhk85);
assign Eugk85 = (Mchk85 & Yg2l85[2]);
assign Mchk85 = (Gi2l85[2] & Tchk85);
assign Tchk85 = (~(Adhk85 & Yg2l85[3]));
assign Adhk85 = (Gi2l85[3] & Hdhk85);
assign Hdhk85 = (~(Odhk85 & Vdhk85));
assign Vdhk85 = (~(Cehk85 & Mb2l85[4]));
assign Cehk85 = (Jehk85 & Z8hk85);
assign Jehk85 = (Ybhk85 | Mb2l85[5]);
assign Odhk85 = (Fchk85 | Mb2l85[7]);
assign Vlgk85 = (Qehk85 & Uogk85);
assign Uogk85 = (~(Yva875 & Xehk85));
assign Xehk85 = (~(Efhk85 & Lfhk85));
assign Qehk85 = (~(M52875 & Wpgk85));
assign M52875 = (!Yva875);
assign Yva875 = (~(Sfhk85 & Zfhk85));
assign Zfhk85 = (~(Gghk85 & Nghk85));
assign Gghk85 = (~(Ughk85 | Kva875));
assign Sfhk85 = (~(Sggk85 & Bhhk85));
assign Bhhk85 = (~(Ihhk85 & Phhk85));
assign Phhk85 = (~(Whhk85 & Dihk85));
assign Dihk85 = (Kihk85 & Lfhk85);
assign Lfhk85 = (~(Rva875 & Rihk85));
assign Kihk85 = (~(Rqgk85 & Yihk85));
assign Whhk85 = (Wpgk85 & Efhk85);
assign Efhk85 = (~(Fjhk85 & Ki9875));
assign Wpgk85 = (Kva875 ? Tjhk85 : Mjhk85);
assign Ihhk85 = (Yihk85 | Rqgk85);
assign Rqgk85 = (Rva875 ? Hkhk85 : Akhk85);
assign Rva875 = (!Ki9875);
assign Yihk85 = (!Yqgk85);
assign Yqgk85 = (Kva875 ? Vkhk85 : Okhk85);
assign Kva875 = (!Ph9875);
assign Ph9875 = (~(Clhk85 & Jlhk85));
assign Jlhk85 = (~(Qlhk85 & Xlhk85));
assign Xlhk85 = (~(Emhk85 & Lmhk85));
assign Lmhk85 = (~(Smhk85 & Tjhk85));
assign Tjhk85 = (Bh9875 ? Mb2l85[18] : Mb2l85[16]);
assign Smhk85 = (~(Mjhk85 | Zmhk85));
assign Zmhk85 = (~(Vkhk85 | Gnhk85));
assign Mjhk85 = (Ih9875 ? Mb2l85[22] : Mb2l85[20]);
assign Emhk85 = (~(Gnhk85 & Vkhk85));
assign Gnhk85 = (!Okhk85);
assign Qlhk85 = (~(Nghk85 & Ih9875));
assign Ih9875 = (!Ughk85);
assign Nghk85 = (~(Yg2l85[11] & Gi2l85[11]));
assign Clhk85 = (~(Bh9875 & Nnhk85));
assign Nnhk85 = (~(Yg2l85[9] & Gi2l85[9]));
assign Vkhk85 = (Bh9875 ? Mb2l85[19] : Mb2l85[17]);
assign Bh9875 = (~(Unhk85 & Yg2l85[8]));
assign Unhk85 = (Gi2l85[8] & Bohk85);
assign Bohk85 = (~(Iohk85 & Yg2l85[9]));
assign Iohk85 = (Gi2l85[9] & Pohk85);
assign Pohk85 = (~(Wohk85 & Dphk85));
assign Dphk85 = (~(Kphk85 & Mb2l85[16]));
assign Kphk85 = (~(Rphk85 | Mb2l85[18]));
assign Rphk85 = (Mb2l85[19] & Yphk85);
assign Wohk85 = (Yphk85 | Mb2l85[19]);
assign Okhk85 = (Ughk85 ? Mb2l85[21] : Mb2l85[23]);
assign Ughk85 = (Fqhk85 & Yg2l85[10]);
assign Fqhk85 = (Gi2l85[10] & Mqhk85);
assign Mqhk85 = (~(Tqhk85 & Yg2l85[11]));
assign Tqhk85 = (Gi2l85[11] & Arhk85);
assign Arhk85 = (~(Hrhk85 & Orhk85));
assign Orhk85 = (~(Vrhk85 & Mb2l85[20]));
assign Vrhk85 = (~(Cshk85 | Mb2l85[22]));
assign Cshk85 = (~(Jshk85 | Mb2l85[21]));
assign Hrhk85 = (~(Mb2l85[21] & Jshk85));
assign Sggk85 = (~(Qshk85 & Xshk85));
assign Qshk85 = (Di9875 & Ki9875);
assign Ki9875 = (~(Ethk85 & Lthk85));
assign Lthk85 = (~(Sthk85 & Zthk85));
assign Zthk85 = (~(Guhk85 & Nuhk85));
assign Nuhk85 = (~(Uuhk85 & Rihk85));
assign Rihk85 = (Wh9875 ? Mb2l85[26] : Mb2l85[24]);
assign Uuhk85 = (~(Fjhk85 | Bvhk85));
assign Bvhk85 = (Akhk85 & Ivhk85);
assign Fjhk85 = (Di9875 ? Mb2l85[30] : Mb2l85[28]);
assign Guhk85 = (Ivhk85 | Akhk85);
assign Akhk85 = (Di9875 ? Mb2l85[31] : Mb2l85[29]);
assign Ivhk85 = (!Hkhk85);
assign Hkhk85 = (Wh9875 ? Mb2l85[27] : Mb2l85[25]);
assign Sthk85 = (~(Xshk85 & Di9875));
assign Xshk85 = (~(Yg2l85[15] & Gi2l85[15]));
assign Ethk85 = (~(Wh9875 & Pvhk85));
assign Pvhk85 = (~(Yg2l85[13] & Gi2l85[13]));
assign Wh9875 = (~(Wvhk85 & Yg2l85[12]));
assign Wvhk85 = (Gi2l85[12] & Dwhk85);
assign Dwhk85 = (~(Kwhk85 & Yg2l85[13]));
assign Kwhk85 = (Gi2l85[13] & Rwhk85);
assign Rwhk85 = (~(Ywhk85 & Fxhk85));
assign Fxhk85 = (~(Mxhk85 & Mb2l85[24]));
assign Mxhk85 = (~(Txhk85 | Mb2l85[26]));
assign Txhk85 = (~(Ayhk85 | Mb2l85[25]));
assign Ywhk85 = (~(Mb2l85[25] & Ayhk85));
assign Di9875 = (~(Hyhk85 & Yg2l85[14]));
assign Hyhk85 = (Gi2l85[14] & Oyhk85);
assign Oyhk85 = (~(Vyhk85 & Yg2l85[15]));
assign Vyhk85 = (Gi2l85[15] & Czhk85);
assign Czhk85 = (~(Jzhk85 & Qzhk85));
assign Qzhk85 = (~(Xzhk85 & Mb2l85[28]));
assign Xzhk85 = (~(E0ik85 | Mb2l85[30]));
assign E0ik85 = (~(L0ik85 | Mb2l85[29]));
assign Jzhk85 = (~(Mb2l85[29] & L0ik85));
assign Hegk85 = (S0ik85 | Z0ik85);
assign Z0ik85 = (T52875 & G1ik85);
assign T52875 = (Ql9875 & Hxa875);
assign S0ik85 = (Ql9875 ? U1ik85 : N1ik85);
assign U1ik85 = (Lm9875 & B2ik85);
assign Uhgk85 = (~(A62875 & Qfgk85));
assign A62875 = (Kjgk85 & Wo9875);
assign Kjgk85 = (!Ql9875);
assign Ql9875 = (I2ik85 & P2ik85);
assign P2ik85 = (~(W2ik85 & D3ik85));
assign D3ik85 = (~(K3ik85 & R3ik85));
assign R3ik85 = (~(Y3ik85 & F4ik85));
assign F4ik85 = (Hxa875 ? G1ik85 : B2ik85);
assign Y3ik85 = (~(N1ik85 | M4ik85));
assign M4ik85 = (Djgk85 & T4ik85);
assign N1ik85 = (Wo9875 ? H5ik85 : A5ik85);
assign K3ik85 = (T4ik85 | Djgk85);
assign Djgk85 = (Wo9875 ? V5ik85 : O5ik85);
assign T4ik85 = (!Wigk85);
assign Wigk85 = (Lm9875 ? J6ik85 : C6ik85);
assign W2ik85 = (~(Qfgk85 & Wo9875));
assign Wo9875 = (~(Q6ik85 & X6ik85));
assign X6ik85 = (~(E7ik85 & L7ik85));
assign E7ik85 = (~(S7ik85 | Vxa875));
assign Q6ik85 = (Qfgk85 | Z7ik85);
assign Z7ik85 = (G8ik85 & N8ik85);
assign N8ik85 = (U8ik85 | H5ik85);
assign H5ik85 = (Rp9875 ? I9ik85 : B9ik85);
assign U8ik85 = (~(A5ik85 & P9ik85));
assign P9ik85 = (~(V5ik85 & W9ik85));
assign A5ik85 = (Mq9875 ? Kaik85 : Daik85);
assign G8ik85 = (W9ik85 | V5ik85);
assign V5ik85 = (Rp9875 ? Yaik85 : Raik85);
assign W9ik85 = (!O5ik85);
assign O5ik85 = (Vxa875 ? Mbik85 : Fbik85);
assign Vxa875 = (!Mq9875);
assign Mq9875 = (~(Tbik85 & Acik85));
assign Acik85 = (~(Hcik85 & Ocik85));
assign Ocik85 = (~(Vcik85 & Cdik85));
assign Cdik85 = (~(Jdik85 & Daik85));
assign Daik85 = (Yp9875 ? Mb2l85[50] : Mb2l85[48]);
assign Jdik85 = (~(Kaik85 | Qdik85));
assign Qdik85 = (~(Mbik85 | Xdik85));
assign Kaik85 = (Fq9875 ? Mb2l85[54] : Mb2l85[52]);
assign Vcik85 = (~(Xdik85 & Mbik85));
assign Xdik85 = (!Fbik85);
assign Hcik85 = (~(L7ik85 & Fq9875));
assign Fq9875 = (!S7ik85);
assign L7ik85 = (Pw8875 | Bui775);
assign Bui775 = (!Gi2l85[27]);
assign Tbik85 = (~(Yp9875 & Eeik85));
assign Eeik85 = (Sk4875 | Sli775);
assign Sli775 = (!Gi2l85[25]);
assign Mbik85 = (Yp9875 ? Mb2l85[51] : Mb2l85[49]);
assign Yp9875 = (~(Leik85 & Yg2l85[24]));
assign Leik85 = (Gi2l85[24] & Seik85);
assign Seik85 = (Zeik85 | Sk4875);
assign Sk4875 = (!Yg2l85[25]);
assign Zeik85 = (~(Gi2l85[25] & Gfik85));
assign Gfik85 = (~(Nfik85 & Ufik85));
assign Ufik85 = (~(Bgik85 & Mb2l85[48]));
assign Bgik85 = (~(Igik85 | Mb2l85[50]));
assign Igik85 = (~(Pgik85 | Mb2l85[49]));
assign Nfik85 = (~(Mb2l85[49] & Pgik85));
assign Fbik85 = (S7ik85 ? Mb2l85[53] : Mb2l85[55]);
assign S7ik85 = (Wgik85 & Yg2l85[26]);
assign Wgik85 = (Gi2l85[26] & Dhik85);
assign Dhik85 = (Khik85 | Pw8875);
assign Pw8875 = (!Yg2l85[27]);
assign Khik85 = (~(Gi2l85[27] & Rhik85));
assign Rhik85 = (~(Yhik85 & Fiik85));
assign Fiik85 = (~(Miik85 & Mb2l85[52]));
assign Miik85 = (~(Tiik85 | Mb2l85[54]));
assign Tiik85 = (~(Ajik85 | Mb2l85[53]));
assign Yhik85 = (~(Mb2l85[53] & Ajik85));
assign I2ik85 = (~(Hjik85 & Ojik85));
assign Ojik85 = (~(Lm9875 | Vjik85));
assign Lm9875 = (!Hxa875);
assign Hxa875 = (~(Ckik85 & Jkik85));
assign Jkik85 = (~(Qkik85 & Xkik85));
assign Xkik85 = (J6ik85 | Elik85);
assign Qkik85 = (Llik85 & Slik85);
assign Slik85 = (~(Zlik85 & Un9875));
assign Zlik85 = (~(Gmik85 | Vjik85));
assign Llik85 = (~(Nmik85 & Umik85));
assign Umik85 = (~(Elik85 & J6ik85));
assign J6ik85 = (Oxa875 ? Inik85 : Bnik85);
assign Elik85 = (!C6ik85);
assign C6ik85 = (Vjik85 ? Wnik85 : Pnik85);
assign Vjik85 = (!Bo9875);
assign Wnik85 = (!Doik85);
assign Nmik85 = (~(Koik85 & B2ik85));
assign B2ik85 = (Oxa875 ? Yoik85 : Roik85);
assign Koik85 = (!G1ik85);
assign G1ik85 = (Bo9875 ? Mpik85 : Fpik85);
assign Bo9875 = (~(Tpik85 & Aqik85));
assign Aqik85 = (~(Hqik85 & Oqik85));
assign Oqik85 = (~(Vqik85 & Crik85));
assign Crik85 = (Jrik85 | Qrik85);
assign Qrik85 = (Un9875 ? Mb2l85[46] : Mb2l85[44]);
assign Un9875 = (!Xrik85);
assign Jrik85 = (~(Fpik85 & Esik85));
assign Esik85 = (~(Pnik85 & Doik85));
assign Vqik85 = (Doik85 | Pnik85);
assign Pnik85 = (Xrik85 ? Mb2l85[45] : Mb2l85[47]);
assign Doik85 = (Nn9875 ? Ssik85 : Lsik85);
assign Hqik85 = (Xrik85 | Gmik85);
assign Tpik85 = (~(Nn9875 & Zsik85));
assign Zsik85 = (~(Yg2l85[21] & Gi2l85[21]));
assign Mpik85 = (Xrik85 ? Mb2l85[44] : Mb2l85[46]);
assign Fpik85 = (Nn9875 ? Mb2l85[42] : Mb2l85[40]);
assign Nn9875 = (~(Gtik85 & Yg2l85[20]));
assign Gtik85 = (Gi2l85[20] & Ntik85);
assign Ntik85 = (~(Utik85 & Yg2l85[21]));
assign Utik85 = (Gi2l85[21] & Buik85);
assign Buik85 = (~(Iuik85 & Puik85));
assign Puik85 = (~(Wuik85 & Mb2l85[40]));
assign Wuik85 = (Dvik85 & Kvik85);
assign Dvik85 = (Ssik85 | Mb2l85[41]);
assign Iuik85 = (Lsik85 | Mb2l85[43]);
assign Ckik85 = (~(Rvik85 & Yvik85));
assign Rvik85 = (~(Fwik85 | Oxa875));
assign Oxa875 = (!Gn9875);
assign Gn9875 = (~(Mwik85 & Twik85));
assign Twik85 = (~(Axik85 & Hxik85));
assign Hxik85 = (~(Oxik85 & Vxik85));
assign Vxik85 = (~(Cyik85 & Yoik85));
assign Yoik85 = (Sm9875 ? Mb2l85[34] : Mb2l85[32]);
assign Cyik85 = (~(Roik85 | Jyik85));
assign Jyik85 = (~(Qyik85 | Inik85));
assign Roik85 = (Zm9875 ? Mb2l85[38] : Mb2l85[36]);
assign Oxik85 = (~(Inik85 & Qyik85));
assign Qyik85 = (!Bnik85);
assign Bnik85 = (Fwik85 ? Mb2l85[37] : Mb2l85[39]);
assign Inik85 = (Sm9875 ? Mb2l85[35] : Mb2l85[33]);
assign Axik85 = (~(Yvik85 & Zm9875));
assign Zm9875 = (!Fwik85);
assign Yvik85 = (~(Yg2l85[19] & Gi2l85[19]));
assign Mwik85 = (~(Sm9875 & Xyik85));
assign Xyik85 = (~(Yg2l85[17] & Gi2l85[17]));
assign Sm9875 = (~(Ezik85 & Yg2l85[16]));
assign Ezik85 = (Gi2l85[16] & Lzik85);
assign Lzik85 = (~(Szik85 & Yg2l85[17]));
assign Szik85 = (Gi2l85[17] & Zzik85);
assign Zzik85 = (~(G0jk85 & N0jk85));
assign N0jk85 = (~(U0jk85 & Mb2l85[32]));
assign U0jk85 = (~(B1jk85 | Mb2l85[34]));
assign B1jk85 = (~(I1jk85 | Mb2l85[33]));
assign G0jk85 = (~(Mb2l85[33] & I1jk85));
assign Fwik85 = (P1jk85 & Yg2l85[18]);
assign P1jk85 = (Gi2l85[18] & W1jk85);
assign W1jk85 = (~(D2jk85 & Yg2l85[19]));
assign D2jk85 = (Gi2l85[19] & K2jk85);
assign K2jk85 = (~(R2jk85 & Y2jk85));
assign Y2jk85 = (~(F3jk85 & Mb2l85[36]));
assign F3jk85 = (~(M3jk85 | Mb2l85[38]));
assign M3jk85 = (~(T3jk85 | Mb2l85[37]));
assign R2jk85 = (~(Mb2l85[37] & T3jk85));
assign Hjik85 = (~(Xrik85 | Gmik85));
assign Xrik85 = (A4jk85 & Yg2l85[22]);
assign A4jk85 = (Gi2l85[22] & H4jk85);
assign H4jk85 = (~(Gmik85 & O4jk85));
assign O4jk85 = (~(V4jk85 & C5jk85));
assign C5jk85 = (~(J5jk85 & Mb2l85[44]));
assign J5jk85 = (~(Q5jk85 | Mb2l85[46]));
assign Q5jk85 = (~(X5jk85 | Mb2l85[45]));
assign V4jk85 = (~(Mb2l85[45] & X5jk85));
assign Gmik85 = (Yg2l85[23] & Gi2l85[23]);
assign Qfgk85 = (E6jk85 & L6jk85);
assign E6jk85 = (Kp9875 & Rp9875);
assign Rp9875 = (~(S6jk85 & Z6jk85));
assign Z6jk85 = (~(G7jk85 & N7jk85));
assign N7jk85 = (~(U7jk85 & B8jk85));
assign B8jk85 = (~(I8jk85 & B9ik85));
assign B9ik85 = (Dp9875 ? Mb2l85[58] : Mb2l85[56]);
assign I8jk85 = (~(I9ik85 | P8jk85));
assign P8jk85 = (Yaik85 & W8jk85);
assign I9ik85 = (Kp9875 ? Mb2l85[62] : Mb2l85[60]);
assign U7jk85 = (W8jk85 | Yaik85);
assign Yaik85 = (Kp9875 ? Mb2l85[63] : Mb2l85[61]);
assign W8jk85 = (!Raik85);
assign Raik85 = (Dp9875 ? Mb2l85[59] : Mb2l85[57]);
assign G7jk85 = (~(L6jk85 & Kp9875));
assign L6jk85 = (~(Yg2l85[31] & Gi2l85[31]));
assign S6jk85 = (~(Dp9875 & D9jk85));
assign D9jk85 = (Geb875 | Xyi775);
assign Xyi775 = (!Gi2l85[29]);
assign Dp9875 = (~(K9jk85 & Yg2l85[28]));
assign K9jk85 = (Gi2l85[28] & R9jk85);
assign R9jk85 = (Y9jk85 | Geb875);
assign Geb875 = (!Yg2l85[29]);
assign Y9jk85 = (~(Gi2l85[29] & Fajk85));
assign Fajk85 = (~(Majk85 & Tajk85));
assign Tajk85 = (~(Abjk85 & Mb2l85[56]));
assign Abjk85 = (~(Hbjk85 | Mb2l85[58]));
assign Hbjk85 = (~(Objk85 | Mb2l85[57]));
assign Majk85 = (~(Mb2l85[57] & Objk85));
assign Kp9875 = (~(Vbjk85 & Yg2l85[30]));
assign Vbjk85 = (Gi2l85[30] & Ccjk85);
assign Ccjk85 = (~(Jcjk85 & Yg2l85[31]));
assign Jcjk85 = (Gi2l85[31] & Qcjk85);
assign Qcjk85 = (~(Xcjk85 & Edjk85));
assign Edjk85 = (~(Ldjk85 & Mb2l85[60]));
assign Ldjk85 = (~(Sdjk85 | Mb2l85[62]));
assign Sdjk85 = (~(Zdjk85 | Mb2l85[61]));
assign Xcjk85 = (~(Mb2l85[61] & Zdjk85));
assign Tse875 = (~(Gejk85 | Ceh775));
assign Ceh775 = (!Vbx775);
assign Gejk85 = (Bj1775 ? vis_primask_o : Ni1775);
assign Bj1775 = (Nejk85 & Uejk85);
assign Uejk85 = (~(Bfjk85 & Ifjk85));
assign Ifjk85 = (N0p675 & Kkf775);
assign Kkf775 = (~(Pfjk85 & Wfjk85));
assign Wfjk85 = (Dgjk85 & Kgjk85);
assign Kgjk85 = (Rgjk85 | Jnf775);
assign Jnf775 = (Ygjk85 & Fhjk85);
assign Fhjk85 = (~(Mhjk85 & Thjk85));
assign Thjk85 = (~(Bvh675 | Rto675));
assign Mhjk85 = (~(Me1775 | Yaw775));
assign Ygjk85 = (X91775 & Aijk85);
assign Aijk85 = (~(Hijk85 & Avy775));
assign Avy775 = (~(D1z675 | Q91775));
assign Hijk85 = (Fvq775 & Gwf775);
assign X91775 = (!Oijk85);
assign Dgjk85 = (Vijk85 | Xnf775);
assign Xnf775 = (Cjjk85 & Jjjk85);
assign Jjjk85 = (Qjjk85 & Xjjk85);
assign Xjjk85 = (~(Z4s775 | Jlv775));
assign Z4s775 = (~(Veg775 | Zry675));
assign Qjjk85 = (Ekjk85 & Xas775);
assign Xas775 = (~(Lkjk85 & Z8a775));
assign Lkjk85 = (~(Me1775 | E5z675));
assign Me1775 = (!Zfa775);
assign Ekjk85 = (~(Skjk85 & O4p675));
assign Skjk85 = (Vxo675 & Zkjk85);
assign Zkjk85 = (~(Gljk85 & K7s775));
assign Gljk85 = (X5p675 | N0p675);
assign Cjjk85 = (Nljk85 & Uljk85);
assign Uljk85 = (~(M3x775 | Bmjk85));
assign Bmjk85 = (Pxf775 & Jf9775);
assign Pxf775 = (Q91775 & Y1z675);
assign M3x775 = (Uag775 & U50775);
assign Nljk85 = (Imjk85 & Pmjk85);
assign Pmjk85 = (~(Zfa775 & U50775));
assign Imjk85 = (N0p675 ? Dnjk85 : Wmjk85);
assign Dnjk85 = (Y1z675 | Q91775);
assign Wmjk85 = (Bbg775 | F3p675);
assign Pfjk85 = (Fsf775 & Knjk85);
assign Knjk85 = (B49775 | Hmf775);
assign Hmf775 = (Rnjk85 & Ynjk85);
assign Ynjk85 = (Mch775 & Fojk85);
assign Fojk85 = (~(Bvh675 & Mojk85));
assign Mojk85 = (~(Tojk85 & Rd1775));
assign Rd1775 = (L2g775 | Mwo675);
assign L2g775 = (!F6g775);
assign Tojk85 = (Apjk85 & Hpjk85);
assign Hpjk85 = (~(Xxq775 & F3p675));
assign Apjk85 = (Wxf775 | D1z675);
assign Wxf775 = (!Zrj775);
assign Mch775 = (~(Opjk85 & Ub1775));
assign Opjk85 = (~(Bbg775 | F3p675));
assign Rnjk85 = (Vpjk85 & Gcl775);
assign Gcl775 = (Ryf775 | Veg775);
assign Vpjk85 = (~(Cqjk85 & Zck775));
assign Cqjk85 = (~(Pw9775 | K1z675));
assign B49775 = (!R2j675);
assign Fsf775 = (N50775 & Jqjk85);
assign Jqjk85 = (~(Qqjk85 & F3p675));
assign Qqjk85 = (Kny675 & Cm2775);
assign N50775 = (!Xqjk85);
assign Bfjk85 = (Tdg775 & Xxq775);
assign Nejk85 = (~(Erjk85 & Xwi675));
assign Erjk85 = (Inb775 & X0a775);
assign X0a775 = (!Pui675);
assign Ni1775 = (~(Lrjk85 & Srjk85));
assign Srjk85 = (~(Zrjk85 & Tdg775));
assign Zrjk85 = (Xxq775 & E0i675);
assign Lrjk85 = (~(Inb775 & Pgp775));
assign Inb775 = (~(Gsjk85 & Nsjk85));
assign Nsjk85 = (~(Usjk85 & F6g775));
assign Usjk85 = (Lsw775 & Xza775);
assign Gsjk85 = (Rux775 | Zry675);
assign Abx775 = (Btjk85 & Itjk85);
assign Itjk85 = (~(Cep675 & Vbx775));
assign Btjk85 = (Vpj775 | Erj775);
assign Vpj775 = (!Wcp675);
assign Dgr675 = (~(Wfr675 & Ptjk85));
assign Ptjk85 = (~(Wtjk85 & Dujk85));
assign Dujk85 = (Kujk85 & Rujk85);
assign Rujk85 = (Yujk85 & Fvjk85);
assign Fvjk85 = (Mvjk85 & Nyz675);
assign Nyz675 = (!hwdata_o[31]);
assign Mvjk85 = (~(hwdata_o[29] | hwdata_o[28]));
assign hwdata_o[28] = (~(Tvjk85 & Awjk85));
assign Awjk85 = (Hwjk85 | Dz0775);
assign Dz0775 = (Owjk85 & Vwjk85);
assign Vwjk85 = (Cxjk85 & Jxjk85);
assign Jxjk85 = (Qxjk85 & Xxjk85);
assign Xxjk85 = (~(vis_r11_o[28] & Eyjk85));
assign Qxjk85 = (Lyjk85 & Syjk85);
assign Syjk85 = (~(vis_r10_o[28] & Zyjk85));
assign Lyjk85 = (~(vis_r9_o[28] & Gzjk85));
assign Cxjk85 = (Nzjk85 & Uzjk85);
assign Uzjk85 = (~(Oom675 & B0kk85));
assign Nzjk85 = (~(vis_r12_o[28] & I0kk85));
assign Owjk85 = (P0kk85 & W0kk85);
assign W0kk85 = (D1kk85 & K1kk85);
assign K1kk85 = (~(vis_r14_o[28] & R1kk85));
assign D1kk85 = (Y1kk85 & F2kk85);
assign F2kk85 = (~(vis_psp_o[26] & M2kk85));
assign Y1kk85 = (~(vis_r8_o[28] & T2kk85));
assign P0kk85 = (B8y675 & A3kk85);
assign A3kk85 = (~(vis_msp_o[26] & H3kk85));
assign B8y675 = (O3kk85 & V3kk85);
assign V3kk85 = (C4kk85 & J4kk85);
assign J4kk85 = (Q4kk85 & X4kk85);
assign X4kk85 = (~(vis_r0_o[28] & E5kk85));
assign Q4kk85 = (~(vis_r2_o[28] & L5kk85));
assign C4kk85 = (S5kk85 & Z5kk85);
assign Z5kk85 = (~(vis_r5_o[28] & G6kk85));
assign S5kk85 = (~(vis_r4_o[28] & N6kk85));
assign O3kk85 = (U6kk85 & B7kk85);
assign B7kk85 = (I7kk85 & P7kk85);
assign P7kk85 = (~(vis_r7_o[28] & W7kk85));
assign I7kk85 = (~(vis_r3_o[28] & D8kk85));
assign U6kk85 = (K8kk85 & R8kk85);
assign R8kk85 = (~(vis_r1_o[28] & Y8kk85));
assign K8kk85 = (~(vis_r6_o[28] & F9kk85));
assign Tvjk85 = (M9kk85 & T9kk85);
assign M9kk85 = (Aakk85 | Lie775);
assign hwdata_o[29] = (~(Hakk85 & Oakk85));
assign Oakk85 = (~(Vakk85 & Ft0775));
assign Ft0775 = (~(Cbkk85 & Jbkk85));
assign Jbkk85 = (Qbkk85 & Xbkk85);
assign Xbkk85 = (Eckk85 & Lckk85);
assign Lckk85 = (~(vis_r11_o[29] & Eyjk85));
assign Eckk85 = (Sckk85 & Zckk85);
assign Zckk85 = (~(vis_r9_o[29] & Gzjk85));
assign Sckk85 = (~(Zpm675 & B0kk85));
assign Qbkk85 = (Gdkk85 & Ndkk85);
assign Ndkk85 = (~(vis_r10_o[29] & Zyjk85));
assign Gdkk85 = (~(vis_psp_o[27] & M2kk85));
assign Cbkk85 = (Udkk85 & Bekk85);
assign Bekk85 = (Iekk85 & Pekk85);
assign Pekk85 = (~(vis_r12_o[29] & I0kk85));
assign Iekk85 = (Wekk85 & Dfkk85);
assign Dfkk85 = (~(vis_msp_o[27] & H3kk85));
assign Wekk85 = (~(vis_r14_o[29] & R1kk85));
assign Udkk85 = (U7y675 & Kfkk85);
assign Kfkk85 = (~(vis_r8_o[29] & T2kk85));
assign U7y675 = (Rfkk85 & Yfkk85);
assign Yfkk85 = (Fgkk85 & Mgkk85);
assign Mgkk85 = (Tgkk85 & Ahkk85);
assign Ahkk85 = (~(vis_r2_o[29] & L5kk85));
assign Tgkk85 = (~(vis_r6_o[29] & F9kk85));
assign Fgkk85 = (Hhkk85 & Ohkk85);
assign Ohkk85 = (~(vis_r5_o[29] & G6kk85));
assign Hhkk85 = (~(vis_r4_o[29] & N6kk85));
assign Rfkk85 = (Vhkk85 & Cikk85);
assign Cikk85 = (Jikk85 & Qikk85);
assign Qikk85 = (~(vis_r1_o[29] & Y8kk85));
assign Jikk85 = (~(vis_r0_o[29] & E5kk85));
assign Vhkk85 = (Xikk85 & Ejkk85);
assign Ejkk85 = (~(vis_r3_o[29] & D8kk85));
assign Xikk85 = (~(vis_r7_o[29] & W7kk85));
assign Hakk85 = (Ljkk85 & Sjkk85);
assign Ljkk85 = (Aakk85 | Nce775);
assign Yujk85 = (~(hwdata_o[27] | hwdata_o[30]));
assign Kujk85 = (Zjkk85 & Gkkk85);
assign Gkkk85 = (~(Cz3775 | hwdata_o[25]));
assign Cz3775 = (!hwdata_o[24]);
assign hwdata_o[24] = (~(Nkkk85 & Ukkk85));
assign Ukkk85 = (Blkk85 | Jdb775);
assign Nkkk85 = (Ilkk85 & Plkk85);
assign Plkk85 = (Aakk85 | W5f775);
assign Ilkk85 = (~(Vakk85 & Qpr775));
assign Qpr775 = (~(Wlkk85 & Dmkk85));
assign Dmkk85 = (Kmkk85 & Rmkk85);
assign Rmkk85 = (Ymkk85 & Fnkk85);
assign Fnkk85 = (~(vis_r11_o[24] & Eyjk85));
assign Ymkk85 = (Mnkk85 & Tnkk85);
assign Tnkk85 = (~(vis_r9_o[24] & Gzjk85));
assign Mnkk85 = (~(Wim675 & B0kk85));
assign Kmkk85 = (Aokk85 & Hokk85);
assign Hokk85 = (~(vis_r10_o[24] & Zyjk85));
assign Aokk85 = (~(vis_psp_o[22] & M2kk85));
assign Wlkk85 = (Ookk85 & Vokk85);
assign Vokk85 = (Cpkk85 & Jpkk85);
assign Jpkk85 = (~(vis_r12_o[24] & I0kk85));
assign Cpkk85 = (Qpkk85 & Xpkk85);
assign Xpkk85 = (~(vis_msp_o[22] & H3kk85));
assign Qpkk85 = (~(vis_r14_o[24] & R1kk85));
assign Ookk85 = (D9y675 & Eqkk85);
assign Eqkk85 = (~(vis_r8_o[24] & T2kk85));
assign D9y675 = (Lqkk85 & Sqkk85);
assign Sqkk85 = (Zqkk85 & Grkk85);
assign Grkk85 = (Nrkk85 & Urkk85);
assign Urkk85 = (~(vis_r2_o[24] & L5kk85));
assign Nrkk85 = (~(vis_r6_o[24] & F9kk85));
assign Zqkk85 = (Bskk85 & Iskk85);
assign Iskk85 = (~(vis_r5_o[24] & G6kk85));
assign Bskk85 = (~(vis_r4_o[24] & N6kk85));
assign Lqkk85 = (Pskk85 & Wskk85);
assign Wskk85 = (Dtkk85 & Ktkk85);
assign Ktkk85 = (~(vis_r1_o[24] & Y8kk85));
assign Dtkk85 = (~(vis_r0_o[24] & E5kk85));
assign Pskk85 = (Rtkk85 & Ytkk85);
assign Ytkk85 = (~(vis_r3_o[24] & D8kk85));
assign Rtkk85 = (~(vis_r7_o[24] & W7kk85));
assign Zjkk85 = (~(hwdata_o[18] | Yw3775));
assign Yw3775 = (!hwdata_o[26]);
assign hwdata_o[26] = (~(Fukk85 & Mukk85));
assign Mukk85 = (Hwjk85 | Rgc775);
assign Rgc775 = (Tukk85 & Avkk85);
assign Avkk85 = (Hvkk85 & Ovkk85);
assign Ovkk85 = (Vvkk85 & Cwkk85);
assign Cwkk85 = (~(vis_r11_o[26] & Eyjk85));
assign Vvkk85 = (Jwkk85 & Qwkk85);
assign Qwkk85 = (~(vis_r9_o[26] & Gzjk85));
assign Jwkk85 = (~(Slm675 & B0kk85));
assign Hvkk85 = (Xwkk85 & Exkk85);
assign Exkk85 = (~(vis_r10_o[26] & Zyjk85));
assign Xwkk85 = (~(vis_psp_o[24] & M2kk85));
assign Tukk85 = (Lxkk85 & Sxkk85);
assign Sxkk85 = (Zxkk85 & Gykk85);
assign Gykk85 = (~(vis_r12_o[26] & I0kk85));
assign Zxkk85 = (Nykk85 & Uykk85);
assign Uykk85 = (~(vis_msp_o[24] & H3kk85));
assign Nykk85 = (~(vis_r14_o[26] & R1kk85));
assign Lxkk85 = (P8y675 & Bzkk85);
assign Bzkk85 = (~(vis_r8_o[26] & T2kk85));
assign P8y675 = (Izkk85 & Pzkk85);
assign Pzkk85 = (Wzkk85 & D0lk85);
assign D0lk85 = (K0lk85 & R0lk85);
assign R0lk85 = (~(vis_r2_o[26] & L5kk85));
assign K0lk85 = (~(vis_r6_o[26] & F9kk85));
assign Wzkk85 = (Y0lk85 & F1lk85);
assign F1lk85 = (~(vis_r5_o[26] & G6kk85));
assign Y0lk85 = (~(vis_r4_o[26] & N6kk85));
assign Izkk85 = (M1lk85 & T1lk85);
assign T1lk85 = (A2lk85 & H2lk85);
assign H2lk85 = (~(vis_r1_o[26] & Y8kk85));
assign A2lk85 = (~(vis_r0_o[26] & E5kk85));
assign M1lk85 = (O2lk85 & V2lk85);
assign V2lk85 = (~(vis_r3_o[26] & D8kk85));
assign O2lk85 = (~(vis_r7_o[26] & W7kk85));
assign Fukk85 = (C3lk85 & J3lk85);
assign C3lk85 = (Aakk85 | Avr775);
assign Wtjk85 = (Q3lk85 & X3lk85);
assign X3lk85 = (E4lk85 & L4lk85);
assign L4lk85 = (S4lk85 & Xk4775);
assign Xk4775 = (hwdata_o[2] & Lnh675);
assign S4lk85 = (~(hwdata_o[16] | G14775));
assign E4lk85 = (hwdata_o[21] & hwdata_o[23]);
assign hwdata_o[23] = (!E04775);
assign E04775 = (Vakk85 ? Plr775 : Elp775);
assign Plr775 = (Z4lk85 & G5lk85);
assign G5lk85 = (N5lk85 & U5lk85);
assign U5lk85 = (B6lk85 & I6lk85);
assign I6lk85 = (~(Lhm675 & B0kk85));
assign B6lk85 = (P6lk85 & W6lk85);
assign W6lk85 = (~(vis_psp_o[21] & M2kk85));
assign P6lk85 = (~(vis_msp_o[21] & H3kk85));
assign N5lk85 = (D7lk85 & K7lk85);
assign K7lk85 = (~(vis_r14_o[23] & R1kk85));
assign D7lk85 = (~(vis_r12_o[23] & I0kk85));
assign Z4lk85 = (R7lk85 & Y7lk85);
assign Y7lk85 = (F8lk85 & M8lk85);
assign M8lk85 = (~(vis_r9_o[23] & Gzjk85));
assign F8lk85 = (T8lk85 & A9lk85);
assign A9lk85 = (~(vis_r11_o[23] & Eyjk85));
assign T8lk85 = (~(vis_r10_o[23] & Zyjk85));
assign R7lk85 = (K9y675 & H9lk85);
assign H9lk85 = (~(vis_r8_o[23] & T2kk85));
assign K9y675 = (O9lk85 & V9lk85);
assign V9lk85 = (Calk85 & Jalk85);
assign Jalk85 = (Qalk85 & Xalk85);
assign Xalk85 = (~(vis_r2_o[23] & L5kk85));
assign Qalk85 = (~(vis_r6_o[23] & F9kk85));
assign Calk85 = (Eblk85 & Lblk85);
assign Lblk85 = (~(vis_r5_o[23] & G6kk85));
assign Eblk85 = (~(vis_r4_o[23] & N6kk85));
assign O9lk85 = (Sblk85 & Zblk85);
assign Zblk85 = (Gclk85 & Nclk85);
assign Nclk85 = (~(vis_r1_o[23] & Y8kk85));
assign Gclk85 = (~(vis_r0_o[23] & E5kk85));
assign Sblk85 = (Uclk85 & Bdlk85);
assign Bdlk85 = (~(vis_r3_o[23] & D8kk85));
assign Uclk85 = (~(vis_r7_o[23] & W7kk85));
assign hwdata_o[21] = (Vakk85 ? Hro775 : U7q775);
assign Hro775 = (~(Idlk85 & Pdlk85));
assign Pdlk85 = (Wdlk85 & Delk85);
assign Delk85 = (Kelk85 & Relk85);
assign Relk85 = (~(vis_r11_o[21] & Eyjk85));
assign Kelk85 = (Yelk85 & Fflk85);
assign Fflk85 = (~(vis_r9_o[21] & Gzjk85));
assign Yelk85 = (~(Pem675 & B0kk85));
assign Wdlk85 = (Mflk85 & Tflk85);
assign Tflk85 = (~(vis_r10_o[21] & Zyjk85));
assign Mflk85 = (~(vis_psp_o[19] & M2kk85));
assign Idlk85 = (Aglk85 & Hglk85);
assign Hglk85 = (Oglk85 & Vglk85);
assign Vglk85 = (~(vis_r12_o[21] & I0kk85));
assign Oglk85 = (Chlk85 & Jhlk85);
assign Jhlk85 = (~(vis_msp_o[19] & H3kk85));
assign Chlk85 = (~(vis_r14_o[21] & R1kk85));
assign Aglk85 = (Y9y675 & Qhlk85);
assign Qhlk85 = (~(vis_r8_o[21] & T2kk85));
assign Y9y675 = (Xhlk85 & Eilk85);
assign Eilk85 = (Lilk85 & Silk85);
assign Silk85 = (Zilk85 & Gjlk85);
assign Gjlk85 = (~(vis_r2_o[21] & L5kk85));
assign Zilk85 = (~(vis_r6_o[21] & F9kk85));
assign Lilk85 = (Njlk85 & Ujlk85);
assign Ujlk85 = (~(vis_r5_o[21] & G6kk85));
assign Njlk85 = (~(vis_r4_o[21] & N6kk85));
assign Xhlk85 = (Bklk85 & Iklk85);
assign Iklk85 = (Pklk85 & Wklk85);
assign Wklk85 = (~(vis_r1_o[21] & Y8kk85));
assign Pklk85 = (~(vis_r0_o[21] & E5kk85));
assign Bklk85 = (Dllk85 & Kllk85);
assign Kllk85 = (~(vis_r3_o[21] & D8kk85));
assign Dllk85 = (~(vis_r7_o[21] & W7kk85));
assign Q3lk85 = (Rllk85 & Yllk85);
assign Yllk85 = (hwdata_o[19] & hwdata_o[20]);
assign hwdata_o[20] = (Vakk85 ? Rpo775 : Apq775);
assign Rpo775 = (~(Fmlk85 & Mmlk85));
assign Mmlk85 = (Tmlk85 & Anlk85);
assign Anlk85 = (Hnlk85 & Onlk85);
assign Onlk85 = (~(vis_r11_o[20] & Eyjk85));
assign Hnlk85 = (Vnlk85 & Colk85);
assign Colk85 = (~(vis_r9_o[20] & Gzjk85));
assign Vnlk85 = (~(Edm675 & B0kk85));
assign Tmlk85 = (Jolk85 & Qolk85);
assign Qolk85 = (~(vis_r10_o[20] & Zyjk85));
assign Jolk85 = (~(vis_psp_o[18] & M2kk85));
assign Fmlk85 = (Xolk85 & Eplk85);
assign Eplk85 = (Lplk85 & Splk85);
assign Splk85 = (~(vis_r12_o[20] & I0kk85));
assign Lplk85 = (Zplk85 & Gqlk85);
assign Gqlk85 = (~(vis_msp_o[18] & H3kk85));
assign Zplk85 = (~(vis_r14_o[20] & R1kk85));
assign Xolk85 = (Fay675 & Nqlk85);
assign Nqlk85 = (~(vis_r8_o[20] & T2kk85));
assign Fay675 = (Uqlk85 & Brlk85);
assign Brlk85 = (Irlk85 & Prlk85);
assign Prlk85 = (Wrlk85 & Dslk85);
assign Dslk85 = (~(vis_r2_o[20] & L5kk85));
assign Wrlk85 = (~(vis_r6_o[20] & F9kk85));
assign Irlk85 = (Kslk85 & Rslk85);
assign Rslk85 = (~(vis_r5_o[20] & G6kk85));
assign Kslk85 = (~(vis_r4_o[20] & N6kk85));
assign Uqlk85 = (Yslk85 & Ftlk85);
assign Ftlk85 = (Mtlk85 & Ttlk85);
assign Ttlk85 = (~(vis_r1_o[20] & Y8kk85));
assign Mtlk85 = (~(vis_r0_o[20] & E5kk85));
assign Yslk85 = (Aulk85 & Hulk85);
assign Hulk85 = (~(vis_r3_o[20] & D8kk85));
assign Aulk85 = (~(vis_r7_o[20] & W7kk85));
assign hwdata_o[19] = (!Oulk85);
assign Oulk85 = (Vakk85 ? Kmd775 : K1d775);
assign Kmd775 = (Vulk85 & Cvlk85);
assign Cvlk85 = (Jvlk85 & Qvlk85);
assign Qvlk85 = (Xvlk85 & Ewlk85);
assign Ewlk85 = (~(vis_r11_o[19] & Eyjk85));
assign Xvlk85 = (Lwlk85 & Swlk85);
assign Swlk85 = (~(vis_r9_o[19] & Gzjk85));
assign Lwlk85 = (~(Tbm675 & B0kk85));
assign Jvlk85 = (Zwlk85 & Gxlk85);
assign Gxlk85 = (~(vis_r10_o[19] & Zyjk85));
assign Zwlk85 = (~(vis_psp_o[17] & M2kk85));
assign Vulk85 = (Nxlk85 & Uxlk85);
assign Uxlk85 = (Bylk85 & Iylk85);
assign Iylk85 = (~(vis_r12_o[19] & I0kk85));
assign Bylk85 = (Pylk85 & Wylk85);
assign Wylk85 = (~(vis_msp_o[17] & H3kk85));
assign Pylk85 = (~(vis_r14_o[19] & R1kk85));
assign Nxlk85 = (Tay675 & Dzlk85);
assign Dzlk85 = (~(vis_r8_o[19] & T2kk85));
assign Tay675 = (Kzlk85 & Rzlk85);
assign Rzlk85 = (Yzlk85 & F0mk85);
assign F0mk85 = (M0mk85 & T0mk85);
assign T0mk85 = (~(vis_r2_o[19] & L5kk85));
assign M0mk85 = (~(vis_r6_o[19] & F9kk85));
assign Yzlk85 = (A1mk85 & H1mk85);
assign H1mk85 = (~(vis_r5_o[19] & G6kk85));
assign A1mk85 = (~(vis_r4_o[19] & N6kk85));
assign Kzlk85 = (O1mk85 & V1mk85);
assign V1mk85 = (C2mk85 & J2mk85);
assign J2mk85 = (~(vis_r1_o[19] & Y8kk85));
assign C2mk85 = (~(vis_r0_o[19] & E5kk85));
assign O1mk85 = (Q2mk85 & X2mk85);
assign X2mk85 = (~(vis_r3_o[19] & D8kk85));
assign Q2mk85 = (~(vis_r7_o[19] & W7kk85));
assign Rllk85 = (~(C64775 | N04875));
assign N04875 = (~(E3mk85 & Zpd875));
assign Zpd875 = (!Ird875);
assign Ird875 = (~(Ycr675 & Ker675));
assign E3mk85 = (Nm4775 & Aar675);
assign Nm4775 = (~(O8r675 | Mbr675));
assign C64775 = (Hwjk85 ? L0p775 : Jwd775);
assign Jwd775 = (!Yap775);
assign Yap775 = (~(L3mk85 & S3mk85));
assign S3mk85 = (Z3mk85 & G4mk85);
assign G4mk85 = (N4mk85 & U4mk85);
assign U4mk85 = (~(vis_r11_o[17] & Eyjk85));
assign N4mk85 = (B5mk85 & I5mk85);
assign I5mk85 = (~(vis_r9_o[17] & Gzjk85));
assign B5mk85 = (~(X8m675 & B0kk85));
assign Z3mk85 = (P5mk85 & W5mk85);
assign W5mk85 = (~(vis_r10_o[17] & Zyjk85));
assign P5mk85 = (~(vis_psp_o[15] & M2kk85));
assign L3mk85 = (D6mk85 & K6mk85);
assign K6mk85 = (R6mk85 & Y6mk85);
assign Y6mk85 = (~(vis_r12_o[17] & I0kk85));
assign R6mk85 = (F7mk85 & M7mk85);
assign M7mk85 = (~(vis_msp_o[15] & H3kk85));
assign F7mk85 = (~(vis_r14_o[17] & R1kk85));
assign D6mk85 = (Hby675 & T7mk85);
assign T7mk85 = (~(vis_r8_o[17] & T2kk85));
assign Hby675 = (A8mk85 & H8mk85);
assign H8mk85 = (O8mk85 & V8mk85);
assign V8mk85 = (C9mk85 & J9mk85);
assign J9mk85 = (~(vis_r2_o[17] & L5kk85));
assign C9mk85 = (~(vis_r6_o[17] & F9kk85));
assign O8mk85 = (Q9mk85 & X9mk85);
assign X9mk85 = (~(vis_r5_o[17] & G6kk85));
assign Q9mk85 = (~(vis_r4_o[17] & N6kk85));
assign A8mk85 = (Eamk85 & Lamk85);
assign Lamk85 = (Samk85 & Zamk85);
assign Zamk85 = (~(vis_r1_o[17] & Y8kk85));
assign Samk85 = (~(vis_r0_o[17] & E5kk85));
assign Eamk85 = (Gbmk85 & Nbmk85);
assign Nbmk85 = (~(vis_r3_o[17] & D8kk85));
assign Gbmk85 = (~(vis_r7_o[17] & W7kk85));
assign hwdata_o[9] = (Ubmk85 ? Rob775 : Z5r775);
assign hwdata_o[8] = (!Gf4775);
assign Gf4775 = (Ubmk85 ? Jdb775 : W5f775);
assign Jdb775 = (!Pgp775);
assign W5f775 = (!Cdp775);
assign Cdp775 = (~(Bcmk85 & Icmk85));
assign Icmk85 = (Pcmk85 & Wcmk85);
assign Wcmk85 = (Ddmk85 & Kdmk85);
assign Kdmk85 = (~(vis_r11_o[8] & Eyjk85));
assign Ddmk85 = (Rdmk85 & Ydmk85);
assign Ydmk85 = (~(vis_r10_o[8] & Zyjk85));
assign Rdmk85 = (~(vis_r9_o[8] & Gzjk85));
assign Pcmk85 = (Femk85 & Memk85);
assign Memk85 = (~(Ewl675 & B0kk85));
assign Femk85 = (~(vis_r12_o[8] & I0kk85));
assign Bcmk85 = (Temk85 & Afmk85);
assign Afmk85 = (Hfmk85 & Ofmk85);
assign Ofmk85 = (~(vis_r14_o[8] & R1kk85));
assign Hfmk85 = (Vfmk85 & Cgmk85);
assign Cgmk85 = (~(vis_psp_o[6] & M2kk85));
assign Vfmk85 = (~(vis_r8_o[8] & T2kk85));
assign Temk85 = (J5y675 & Jgmk85);
assign Jgmk85 = (~(vis_msp_o[6] & H3kk85));
assign J5y675 = (Qgmk85 & Xgmk85);
assign Xgmk85 = (Ehmk85 & Lhmk85);
assign Lhmk85 = (Shmk85 & Zhmk85);
assign Zhmk85 = (~(vis_r0_o[8] & E5kk85));
assign Shmk85 = (~(vis_r2_o[8] & L5kk85));
assign Ehmk85 = (Gimk85 & Nimk85);
assign Nimk85 = (~(vis_r5_o[8] & G6kk85));
assign Gimk85 = (~(vis_r4_o[8] & N6kk85));
assign Qgmk85 = (Uimk85 & Bjmk85);
assign Bjmk85 = (Ijmk85 & Pjmk85);
assign Pjmk85 = (~(vis_r7_o[8] & W7kk85));
assign Ijmk85 = (~(vis_r3_o[8] & D8kk85));
assign Uimk85 = (Wjmk85 & Dkmk85);
assign Dkmk85 = (~(vis_r1_o[8] & Y8kk85));
assign Wjmk85 = (~(vis_r6_o[8] & F9kk85));
assign hwdata_o[7] = (Oxh675 & Ajp775);
assign hwdata_o[6] = (Oxh675 & Zep775);
assign hwdata_o[5] = (Oxh675 & U7q775);
assign hwdata_o[4] = (Oxh675 & Apq775);
assign hwdata_o[3] = (Oxh675 & Fbp775);
assign hwdata_o[31] = (~(Kkmk85 & Rkmk85));
assign Rkmk85 = (Blkk85 | Elp775);
assign Kkmk85 = (Ykmk85 & Flmk85);
assign Flmk85 = (~(Vakk85 & Pig775));
assign Pig775 = (~(Mlmk85 & Tlmk85));
assign Tlmk85 = (Ammk85 & Hmmk85);
assign Hmmk85 = (Ommk85 & Vmmk85);
assign Vmmk85 = (~(vis_r11_o[31] & Eyjk85));
assign Ommk85 = (Cnmk85 & Jnmk85);
assign Jnmk85 = (~(vis_r10_o[31] & Zyjk85));
assign Cnmk85 = (~(vis_r9_o[31] & Gzjk85));
assign Ammk85 = (Qnmk85 & Xnmk85);
assign Xnmk85 = (~(Vsm675 & B0kk85));
assign Qnmk85 = (~(vis_r12_o[31] & I0kk85));
assign Mlmk85 = (Eomk85 & Lomk85);
assign Lomk85 = (Somk85 & Zomk85);
assign Zomk85 = (~(vis_r14_o[31] & R1kk85));
assign Somk85 = (Gpmk85 & Npmk85);
assign Npmk85 = (~(vis_psp_o[29] & M2kk85));
assign Gpmk85 = (~(vis_r8_o[31] & T2kk85));
assign Eomk85 = (Z6y675 & Upmk85);
assign Upmk85 = (~(vis_msp_o[29] & H3kk85));
assign Z6y675 = (Bqmk85 & Iqmk85);
assign Iqmk85 = (Pqmk85 & Wqmk85);
assign Wqmk85 = (Drmk85 & Krmk85);
assign Krmk85 = (~(vis_r0_o[31] & E5kk85));
assign Drmk85 = (~(vis_r2_o[31] & L5kk85));
assign Pqmk85 = (Rrmk85 & Yrmk85);
assign Yrmk85 = (~(vis_r5_o[31] & G6kk85));
assign Rrmk85 = (~(vis_r4_o[31] & N6kk85));
assign Bqmk85 = (Fsmk85 & Msmk85);
assign Msmk85 = (Tsmk85 & Atmk85);
assign Atmk85 = (~(vis_r7_o[31] & W7kk85));
assign Tsmk85 = (~(vis_r3_o[31] & D8kk85));
assign Fsmk85 = (Htmk85 & Otmk85);
assign Otmk85 = (~(vis_r1_o[31] & Y8kk85));
assign Htmk85 = (~(vis_r6_o[31] & F9kk85));
assign Ykmk85 = (Aakk85 | Saf775);
assign hwdata_o[30] = (~(Vtmk85 & Cumk85));
assign Cumk85 = (Blkk85 | Gsc775);
assign Vtmk85 = (Jumk85 & Qumk85);
assign Qumk85 = (Hwjk85 | Y2c775);
assign Y2c775 = (!Ocp775);
assign Ocp775 = (~(Xumk85 & Evmk85));
assign Evmk85 = (Lvmk85 & Svmk85);
assign Svmk85 = (Zvmk85 & Gwmk85);
assign Gwmk85 = (~(vis_r11_o[30] & Eyjk85));
assign Zvmk85 = (Nwmk85 & Uwmk85);
assign Uwmk85 = (~(vis_r10_o[30] & Zyjk85));
assign Nwmk85 = (~(vis_r9_o[30] & Gzjk85));
assign Lvmk85 = (Bxmk85 & Ixmk85);
assign Ixmk85 = (~(Krm675 & B0kk85));
assign Bxmk85 = (~(vis_r12_o[30] & I0kk85));
assign Xumk85 = (Pxmk85 & Wxmk85);
assign Wxmk85 = (Dymk85 & Kymk85);
assign Kymk85 = (~(vis_r14_o[30] & R1kk85));
assign Dymk85 = (Rymk85 & Yymk85);
assign Yymk85 = (~(vis_psp_o[28] & M2kk85));
assign Rymk85 = (~(vis_r8_o[30] & T2kk85));
assign Pxmk85 = (G7y675 & Fzmk85);
assign Fzmk85 = (~(vis_msp_o[28] & H3kk85));
assign G7y675 = (Mzmk85 & Tzmk85);
assign Tzmk85 = (A0nk85 & H0nk85);
assign H0nk85 = (O0nk85 & V0nk85);
assign V0nk85 = (~(vis_r0_o[30] & E5kk85));
assign O0nk85 = (~(vis_r2_o[30] & L5kk85));
assign A0nk85 = (C1nk85 & J1nk85);
assign J1nk85 = (~(vis_r5_o[30] & G6kk85));
assign C1nk85 = (~(vis_r4_o[30] & N6kk85));
assign Mzmk85 = (Q1nk85 & X1nk85);
assign X1nk85 = (E2nk85 & L2nk85);
assign L2nk85 = (~(vis_r7_o[30] & W7kk85));
assign E2nk85 = (~(vis_r3_o[30] & D8kk85));
assign Q1nk85 = (S2nk85 & Z2nk85);
assign Z2nk85 = (~(vis_r1_o[30] & Y8kk85));
assign S2nk85 = (~(vis_r6_o[30] & F9kk85));
assign Jumk85 = (Aakk85 | K7e775);
assign hwdata_o[2] = (~(Me8775 | Neq775));
assign hwdata_o[27] = (~(G3nk85 & N3nk85));
assign N3nk85 = (Blkk85 | K1d775);
assign G3nk85 = (U3nk85 & B4nk85);
assign B4nk85 = (~(Vakk85 & Cir775));
assign Cir775 = (~(I4nk85 & P4nk85));
assign P4nk85 = (W4nk85 & D5nk85);
assign D5nk85 = (K5nk85 & R5nk85);
assign R5nk85 = (~(vis_r11_o[27] & Eyjk85));
assign K5nk85 = (Y5nk85 & F6nk85);
assign F6nk85 = (~(vis_r9_o[27] & Gzjk85));
assign Y5nk85 = (~(Dnm675 & B0kk85));
assign W4nk85 = (M6nk85 & T6nk85);
assign T6nk85 = (~(vis_r10_o[27] & Zyjk85));
assign M6nk85 = (~(vis_psp_o[25] & M2kk85));
assign I4nk85 = (A7nk85 & H7nk85);
assign H7nk85 = (O7nk85 & V7nk85);
assign V7nk85 = (~(vis_r12_o[27] & I0kk85));
assign O7nk85 = (C8nk85 & J8nk85);
assign J8nk85 = (~(vis_msp_o[25] & H3kk85));
assign C8nk85 = (~(vis_r14_o[27] & R1kk85));
assign A7nk85 = (I8y675 & Q8nk85);
assign Q8nk85 = (~(vis_r8_o[27] & T2kk85));
assign I8y675 = (X8nk85 & E9nk85);
assign E9nk85 = (L9nk85 & S9nk85);
assign S9nk85 = (Z9nk85 & Gank85);
assign Gank85 = (~(vis_r2_o[27] & L5kk85));
assign Z9nk85 = (~(vis_r6_o[27] & F9kk85));
assign L9nk85 = (Nank85 & Uank85);
assign Uank85 = (~(vis_r5_o[27] & G6kk85));
assign Nank85 = (~(vis_r4_o[27] & N6kk85));
assign X8nk85 = (Bbnk85 & Ibnk85);
assign Ibnk85 = (Pbnk85 & Wbnk85);
assign Wbnk85 = (~(vis_r1_o[27] & Y8kk85));
assign Pbnk85 = (~(vis_r0_o[27] & E5kk85));
assign Bbnk85 = (Dcnk85 & Kcnk85);
assign Kcnk85 = (~(vis_r3_o[27] & D8kk85));
assign Dcnk85 = (~(vis_r7_o[27] & W7kk85));
assign U3nk85 = (Aakk85 | Xoe775);
assign hwdata_o[25] = (~(Rcnk85 & Ycnk85));
assign Ycnk85 = (Blkk85 | L0p775);
assign L0p775 = (!Rob775);
assign Rcnk85 = (Fdnk85 & Mdnk85);
assign Mdnk85 = (Hwjk85 | Wmc775);
assign Wmc775 = (!Hcp775);
assign Hcp775 = (~(Tdnk85 & Aenk85));
assign Aenk85 = (Henk85 & Oenk85);
assign Oenk85 = (Venk85 & Cfnk85);
assign Cfnk85 = (~(vis_r11_o[25] & Eyjk85));
assign Venk85 = (Jfnk85 & Qfnk85);
assign Qfnk85 = (~(vis_r9_o[25] & Gzjk85));
assign Jfnk85 = (~(Hkm675 & B0kk85));
assign Henk85 = (Xfnk85 & Egnk85);
assign Egnk85 = (~(vis_r10_o[25] & Zyjk85));
assign Xfnk85 = (~(vis_psp_o[23] & M2kk85));
assign Tdnk85 = (Lgnk85 & Sgnk85);
assign Sgnk85 = (Zgnk85 & Ghnk85);
assign Ghnk85 = (~(vis_r12_o[25] & I0kk85));
assign Zgnk85 = (Nhnk85 & Uhnk85);
assign Uhnk85 = (~(vis_msp_o[23] & H3kk85));
assign Nhnk85 = (~(vis_r14_o[25] & R1kk85));
assign Lgnk85 = (W8y675 & Bink85);
assign Bink85 = (~(vis_r8_o[25] & T2kk85));
assign W8y675 = (Iink85 & Pink85);
assign Pink85 = (Wink85 & Djnk85);
assign Djnk85 = (Kjnk85 & Rjnk85);
assign Rjnk85 = (~(vis_r2_o[25] & L5kk85));
assign Kjnk85 = (~(vis_r6_o[25] & F9kk85));
assign Wink85 = (Yjnk85 & Fknk85);
assign Fknk85 = (~(vis_r5_o[25] & G6kk85));
assign Yjnk85 = (~(vis_r4_o[25] & N6kk85));
assign Iink85 = (Mknk85 & Tknk85);
assign Tknk85 = (Alnk85 & Hlnk85);
assign Hlnk85 = (~(vis_r1_o[25] & Y8kk85));
assign Alnk85 = (~(vis_r0_o[25] & E5kk85));
assign Mknk85 = (Olnk85 & Vlnk85);
assign Vlnk85 = (~(vis_r3_o[25] & D8kk85));
assign Olnk85 = (~(vis_r7_o[25] & W7kk85));
assign Fdnk85 = (~(Cmnk85 & Z5r775));
assign Z5r775 = (~(Jmnk85 & Qmnk85));
assign Qmnk85 = (Xmnk85 & Ennk85);
assign Ennk85 = (Lnnk85 & Snnk85);
assign Snnk85 = (~(Oxl675 & B0kk85));
assign Lnnk85 = (Znnk85 & Gonk85);
assign Gonk85 = (~(vis_psp_o[7] & M2kk85));
assign Znnk85 = (~(vis_msp_o[7] & H3kk85));
assign Xmnk85 = (Nonk85 & Uonk85);
assign Uonk85 = (~(vis_r14_o[9] & R1kk85));
assign Nonk85 = (~(vis_r12_o[9] & I0kk85));
assign Jmnk85 = (Bpnk85 & Ipnk85);
assign Ipnk85 = (Ppnk85 & Wpnk85);
assign Wpnk85 = (~(vis_r9_o[9] & Gzjk85));
assign Ppnk85 = (Dqnk85 & Kqnk85);
assign Kqnk85 = (~(vis_r11_o[9] & Eyjk85));
assign Dqnk85 = (~(vis_r10_o[9] & Zyjk85));
assign Bpnk85 = (V4y675 & Rqnk85);
assign Rqnk85 = (~(vis_r8_o[9] & T2kk85));
assign V4y675 = (Yqnk85 & Frnk85);
assign Frnk85 = (Mrnk85 & Trnk85);
assign Trnk85 = (Asnk85 & Hsnk85);
assign Hsnk85 = (~(vis_r2_o[9] & L5kk85));
assign Asnk85 = (~(vis_r6_o[9] & F9kk85));
assign Mrnk85 = (Osnk85 & Vsnk85);
assign Vsnk85 = (~(vis_r5_o[9] & G6kk85));
assign Osnk85 = (~(vis_r4_o[9] & N6kk85));
assign Yqnk85 = (Ctnk85 & Jtnk85);
assign Jtnk85 = (Qtnk85 & Xtnk85);
assign Xtnk85 = (~(vis_r1_o[9] & Y8kk85));
assign Qtnk85 = (~(vis_r0_o[9] & E5kk85));
assign Ctnk85 = (Eunk85 & Lunk85);
assign Lunk85 = (~(vis_r3_o[9] & D8kk85));
assign Eunk85 = (~(vis_r7_o[9] & W7kk85));
assign Cmnk85 = (!Aakk85);
assign Aakk85 = (~(Sunk85 & Oxh675));
assign hwdata_o[22] = (!G14775);
assign G14775 = (Vakk85 ? P7d775 : Gsc775);
assign P7d775 = (!Vcp775);
assign Vcp775 = (~(Zunk85 & Gvnk85));
assign Gvnk85 = (Nvnk85 & Uvnk85);
assign Uvnk85 = (Bwnk85 & Iwnk85);
assign Iwnk85 = (~(vis_r11_o[22] & Eyjk85));
assign Bwnk85 = (Pwnk85 & Wwnk85);
assign Wwnk85 = (~(vis_r9_o[22] & Gzjk85));
assign Pwnk85 = (~(Agm675 & B0kk85));
assign Nvnk85 = (Dxnk85 & Kxnk85);
assign Kxnk85 = (~(vis_r10_o[22] & Zyjk85));
assign Dxnk85 = (~(vis_psp_o[20] & M2kk85));
assign Zunk85 = (Rxnk85 & Yxnk85);
assign Yxnk85 = (Fynk85 & Mynk85);
assign Mynk85 = (~(vis_r12_o[22] & I0kk85));
assign Fynk85 = (Tynk85 & Aznk85);
assign Aznk85 = (~(vis_msp_o[20] & H3kk85));
assign Tynk85 = (~(vis_r14_o[22] & R1kk85));
assign Rxnk85 = (R9y675 & Hznk85);
assign Hznk85 = (~(vis_r8_o[22] & T2kk85));
assign R9y675 = (Oznk85 & Vznk85);
assign Vznk85 = (C0ok85 & J0ok85);
assign J0ok85 = (Q0ok85 & X0ok85);
assign X0ok85 = (~(vis_r2_o[22] & L5kk85));
assign Q0ok85 = (~(vis_r6_o[22] & F9kk85));
assign C0ok85 = (E1ok85 & L1ok85);
assign L1ok85 = (~(vis_r5_o[22] & G6kk85));
assign E1ok85 = (~(vis_r4_o[22] & N6kk85));
assign Oznk85 = (S1ok85 & Z1ok85);
assign Z1ok85 = (G2ok85 & N2ok85);
assign N2ok85 = (~(vis_r1_o[22] & Y8kk85));
assign G2ok85 = (~(vis_r0_o[22] & E5kk85));
assign S1ok85 = (U2ok85 & B3ok85);
assign B3ok85 = (~(vis_r3_o[22] & D8kk85));
assign U2ok85 = (~(vis_r7_o[22] & W7kk85));
assign hwdata_o[1] = (Oxh675 & Rob775);
assign Rob775 = (~(I3ok85 & P3ok85));
assign P3ok85 = (W3ok85 & D4ok85);
assign D4ok85 = (K4ok85 & R4ok85);
assign R4ok85 = (~(vis_r10_o[1] & Zyjk85));
assign K4ok85 = (~(Mml675 & B0kk85));
assign W3ok85 = (Y4ok85 & F5ok85);
assign F5ok85 = (~(vis_r12_o[1] & I0kk85));
assign Y4ok85 = (~(vis_r11_o[1] & Eyjk85));
assign I3ok85 = (M5ok85 & T5ok85);
assign T5ok85 = (A6ok85 & H6ok85);
assign H6ok85 = (~(vis_r8_o[1] & T2kk85));
assign A6ok85 = (~(vis_r9_o[1] & Gzjk85));
assign M5ok85 = (May675 & O6ok85);
assign O6ok85 = (~(vis_r14_o[1] & R1kk85));
assign May675 = (V6ok85 & C7ok85);
assign C7ok85 = (J7ok85 & Q7ok85);
assign Q7ok85 = (X7ok85 & E8ok85);
assign E8ok85 = (~(vis_r0_o[1] & E5kk85));
assign X7ok85 = (~(vis_r2_o[1] & L5kk85));
assign J7ok85 = (L8ok85 & S8ok85);
assign S8ok85 = (~(vis_r5_o[1] & G6kk85));
assign L8ok85 = (~(vis_r4_o[1] & N6kk85));
assign V6ok85 = (Z8ok85 & G9ok85);
assign G9ok85 = (N9ok85 & U9ok85);
assign U9ok85 = (~(vis_r7_o[1] & W7kk85));
assign N9ok85 = (~(vis_r3_o[1] & D8kk85));
assign Z8ok85 = (Baok85 & Iaok85);
assign Iaok85 = (~(vis_r1_o[1] & Y8kk85));
assign Baok85 = (~(vis_r6_o[1] & F9kk85));
assign hwdata_o[18] = (!A54775);
assign A54775 = (Vakk85 ? Grd775 : Neq775);
assign Grd775 = (!Sep775);
assign Sep775 = (~(Paok85 & Waok85));
assign Waok85 = (Dbok85 & Kbok85);
assign Kbok85 = (Rbok85 & Ybok85);
assign Ybok85 = (~(vis_r11_o[18] & Eyjk85));
assign Rbok85 = (Fcok85 & Mcok85);
assign Mcok85 = (~(vis_r9_o[18] & Gzjk85));
assign Fcok85 = (~(Iam675 & B0kk85));
assign Dbok85 = (Tcok85 & Adok85);
assign Adok85 = (~(vis_r10_o[18] & Zyjk85));
assign Tcok85 = (~(vis_psp_o[16] & M2kk85));
assign Paok85 = (Hdok85 & Odok85);
assign Odok85 = (Vdok85 & Ceok85);
assign Ceok85 = (~(vis_r12_o[18] & I0kk85));
assign Vdok85 = (Jeok85 & Qeok85);
assign Qeok85 = (~(vis_msp_o[16] & H3kk85));
assign Jeok85 = (~(vis_r14_o[18] & R1kk85));
assign Hdok85 = (Aby675 & Xeok85);
assign Xeok85 = (~(vis_r8_o[18] & T2kk85));
assign Aby675 = (Efok85 & Lfok85);
assign Lfok85 = (Sfok85 & Zfok85);
assign Zfok85 = (Ggok85 & Ngok85);
assign Ngok85 = (~(vis_r2_o[18] & L5kk85));
assign Ggok85 = (~(vis_r6_o[18] & F9kk85));
assign Sfok85 = (Ugok85 & Bhok85);
assign Bhok85 = (~(vis_r5_o[18] & G6kk85));
assign Ugok85 = (~(vis_r4_o[18] & N6kk85));
assign Efok85 = (Ihok85 & Phok85);
assign Phok85 = (Whok85 & Diok85);
assign Diok85 = (~(vis_r1_o[18] & Y8kk85));
assign Whok85 = (~(vis_r0_o[18] & E5kk85));
assign Ihok85 = (Kiok85 & Riok85);
assign Riok85 = (~(vis_r3_o[18] & D8kk85));
assign Kiok85 = (~(vis_r7_o[18] & W7kk85));
assign hwdata_o[16] = (Hwjk85 ? Pgp775 : Boo775);
assign Hwjk85 = (!Vakk85);
assign Vakk85 = (~(Me8775 | Yiok85));
assign Boo775 = (~(Fjok85 & Mjok85));
assign Mjok85 = (Tjok85 & Akok85);
assign Akok85 = (Hkok85 & Okok85);
assign Okok85 = (~(vis_r11_o[16] & Eyjk85));
assign Hkok85 = (Vkok85 & Clok85);
assign Clok85 = (~(vis_r9_o[16] & Gzjk85));
assign Vkok85 = (~(M7m675 & B0kk85));
assign Tjok85 = (Jlok85 & Qlok85);
assign Qlok85 = (~(vis_r10_o[16] & Zyjk85));
assign Jlok85 = (~(vis_psp_o[14] & M2kk85));
assign Fjok85 = (Xlok85 & Emok85);
assign Emok85 = (Lmok85 & Smok85);
assign Smok85 = (~(vis_r12_o[16] & I0kk85));
assign Lmok85 = (Zmok85 & Gnok85);
assign Gnok85 = (~(vis_msp_o[14] & H3kk85));
assign Zmok85 = (~(vis_r14_o[16] & R1kk85));
assign Xlok85 = (Oby675 & Nnok85);
assign Nnok85 = (~(vis_r8_o[16] & T2kk85));
assign Oby675 = (Unok85 & Book85);
assign Book85 = (Iook85 & Pook85);
assign Pook85 = (Wook85 & Dpok85);
assign Dpok85 = (~(vis_r2_o[16] & L5kk85));
assign Wook85 = (~(vis_r6_o[16] & F9kk85));
assign Iook85 = (Kpok85 & Rpok85);
assign Rpok85 = (~(vis_r5_o[16] & G6kk85));
assign Kpok85 = (~(vis_r4_o[16] & N6kk85));
assign Unok85 = (Ypok85 & Fqok85);
assign Fqok85 = (Mqok85 & Tqok85);
assign Tqok85 = (~(vis_r1_o[16] & Y8kk85));
assign Mqok85 = (~(vis_r0_o[16] & E5kk85));
assign Ypok85 = (Arok85 & Hrok85);
assign Hrok85 = (~(vis_r3_o[16] & D8kk85));
assign Arok85 = (~(vis_r7_o[16] & W7kk85));
assign hwdata_o[15] = (!Z74775);
assign Z74775 = (Ubmk85 ? Elp775 : Saf775);
assign Elp775 = (!Ajp775);
assign Ajp775 = (~(Orok85 & Vrok85));
assign Vrok85 = (Csok85 & Jsok85);
assign Jsok85 = (Qsok85 & Xsok85);
assign Xsok85 = (~(vis_r11_o[7] & Eyjk85));
assign Qsok85 = (Etok85 & Ltok85);
assign Ltok85 = (~(vis_r9_o[7] & Gzjk85));
assign Etok85 = (~(Uul675 & B0kk85));
assign Csok85 = (Stok85 & Ztok85);
assign Ztok85 = (~(vis_r10_o[7] & Zyjk85));
assign Stok85 = (~(vis_psp_o[5] & M2kk85));
assign Orok85 = (Guok85 & Nuok85);
assign Nuok85 = (Uuok85 & Bvok85);
assign Bvok85 = (~(vis_r12_o[7] & I0kk85));
assign Uuok85 = (Ivok85 & Pvok85);
assign Pvok85 = (~(vis_msp_o[5] & H3kk85));
assign Ivok85 = (~(vis_r14_o[7] & R1kk85));
assign Guok85 = (Q5y675 & Wvok85);
assign Wvok85 = (~(vis_r8_o[7] & T2kk85));
assign Q5y675 = (Dwok85 & Kwok85);
assign Kwok85 = (Rwok85 & Ywok85);
assign Ywok85 = (Fxok85 & Mxok85);
assign Mxok85 = (~(vis_r0_o[7] & E5kk85));
assign Fxok85 = (~(vis_r2_o[7] & L5kk85));
assign Rwok85 = (Txok85 & Ayok85);
assign Ayok85 = (~(vis_r5_o[7] & G6kk85));
assign Txok85 = (~(vis_r4_o[7] & N6kk85));
assign Dwok85 = (Hyok85 & Oyok85);
assign Oyok85 = (Vyok85 & Czok85);
assign Czok85 = (~(vis_r7_o[7] & W7kk85));
assign Vyok85 = (~(vis_r3_o[7] & D8kk85));
assign Hyok85 = (Jzok85 & Qzok85);
assign Qzok85 = (~(vis_r1_o[7] & Y8kk85));
assign Jzok85 = (~(vis_r6_o[7] & F9kk85));
assign Saf775 = (Xzok85 & E0pk85);
assign E0pk85 = (L0pk85 & S0pk85);
assign S0pk85 = (Z0pk85 & G1pk85);
assign G1pk85 = (~(vis_r11_o[15] & Eyjk85));
assign Z0pk85 = (N1pk85 & U1pk85);
assign U1pk85 = (~(vis_r10_o[15] & Zyjk85));
assign N1pk85 = (~(vis_r9_o[15] & Gzjk85));
assign L0pk85 = (B2pk85 & I2pk85);
assign I2pk85 = (~(B6m675 & B0kk85));
assign B2pk85 = (~(vis_r12_o[15] & I0kk85));
assign Xzok85 = (P2pk85 & W2pk85);
assign W2pk85 = (D3pk85 & K3pk85);
assign K3pk85 = (~(vis_r14_o[15] & R1kk85));
assign D3pk85 = (R3pk85 & Y3pk85);
assign Y3pk85 = (~(vis_psp_o[13] & M2kk85));
assign R3pk85 = (~(vis_r8_o[15] & T2kk85));
assign P2pk85 = (Vby675 & F4pk85);
assign F4pk85 = (~(vis_msp_o[13] & H3kk85));
assign Vby675 = (M4pk85 & T4pk85);
assign T4pk85 = (A5pk85 & H5pk85);
assign H5pk85 = (O5pk85 & V5pk85);
assign V5pk85 = (~(vis_r0_o[15] & E5kk85));
assign O5pk85 = (~(vis_r2_o[15] & L5kk85));
assign A5pk85 = (C6pk85 & J6pk85);
assign J6pk85 = (~(vis_r5_o[15] & G6kk85));
assign C6pk85 = (~(vis_r4_o[15] & N6kk85));
assign M4pk85 = (Q6pk85 & X6pk85);
assign X6pk85 = (E7pk85 & L7pk85);
assign L7pk85 = (~(vis_r7_o[15] & W7kk85));
assign E7pk85 = (~(vis_r3_o[15] & D8kk85));
assign Q6pk85 = (S7pk85 & Z7pk85);
assign Z7pk85 = (~(vis_r1_o[15] & Y8kk85));
assign S7pk85 = (~(vis_r6_o[15] & F9kk85));
assign hwdata_o[14] = (!B94775);
assign B94775 = (Ubmk85 ? Gsc775 : K7e775);
assign Gsc775 = (!Zep775);
assign Zep775 = (~(G8pk85 & N8pk85));
assign N8pk85 = (U8pk85 & B9pk85);
assign B9pk85 = (I9pk85 & P9pk85);
assign P9pk85 = (~(vis_r11_o[6] & Eyjk85));
assign I9pk85 = (W9pk85 & Dapk85);
assign Dapk85 = (~(vis_r9_o[6] & Gzjk85));
assign W9pk85 = (~(Ktl675 & B0kk85));
assign U8pk85 = (Kapk85 & Rapk85);
assign Rapk85 = (~(vis_r10_o[6] & Zyjk85));
assign Kapk85 = (~(vis_psp_o[4] & M2kk85));
assign G8pk85 = (Yapk85 & Fbpk85);
assign Fbpk85 = (Mbpk85 & Tbpk85);
assign Tbpk85 = (~(vis_r12_o[6] & I0kk85));
assign Mbpk85 = (Acpk85 & Hcpk85);
assign Hcpk85 = (~(vis_msp_o[4] & H3kk85));
assign Acpk85 = (~(vis_r14_o[6] & R1kk85));
assign Yapk85 = (X5y675 & Ocpk85);
assign Ocpk85 = (~(vis_r8_o[6] & T2kk85));
assign X5y675 = (Vcpk85 & Cdpk85);
assign Cdpk85 = (Jdpk85 & Qdpk85);
assign Qdpk85 = (Xdpk85 & Eepk85);
assign Eepk85 = (~(vis_r0_o[6] & E5kk85));
assign Xdpk85 = (~(vis_r2_o[6] & L5kk85));
assign Jdpk85 = (Lepk85 & Sepk85);
assign Sepk85 = (~(vis_r5_o[6] & G6kk85));
assign Lepk85 = (~(vis_r4_o[6] & N6kk85));
assign Vcpk85 = (Zepk85 & Gfpk85);
assign Gfpk85 = (Nfpk85 & Ufpk85);
assign Ufpk85 = (~(vis_r7_o[6] & W7kk85));
assign Nfpk85 = (~(vis_r3_o[6] & D8kk85));
assign Zepk85 = (Bgpk85 & Igpk85);
assign Igpk85 = (~(vis_r1_o[6] & Y8kk85));
assign Bgpk85 = (~(vis_r6_o[6] & F9kk85));
assign K7e775 = (!Gfp775);
assign Gfp775 = (~(Pgpk85 & Wgpk85));
assign Wgpk85 = (Dhpk85 & Khpk85);
assign Khpk85 = (Rhpk85 & Yhpk85);
assign Yhpk85 = (~(vis_r11_o[14] & Eyjk85));
assign Rhpk85 = (Fipk85 & Mipk85);
assign Mipk85 = (~(vis_r10_o[14] & Zyjk85));
assign Fipk85 = (~(vis_r9_o[14] & Gzjk85));
assign Dhpk85 = (Tipk85 & Ajpk85);
assign Ajpk85 = (~(Q4m675 & B0kk85));
assign Tipk85 = (~(vis_r12_o[14] & I0kk85));
assign Pgpk85 = (Hjpk85 & Ojpk85);
assign Ojpk85 = (Vjpk85 & Ckpk85);
assign Ckpk85 = (~(vis_r14_o[14] & R1kk85));
assign Vjpk85 = (Jkpk85 & Qkpk85);
assign Qkpk85 = (~(vis_psp_o[12] & M2kk85));
assign Jkpk85 = (~(vis_r8_o[14] & T2kk85));
assign Hjpk85 = (Ccy675 & Xkpk85);
assign Xkpk85 = (~(vis_msp_o[12] & H3kk85));
assign Ccy675 = (Elpk85 & Llpk85);
assign Llpk85 = (Slpk85 & Zlpk85);
assign Zlpk85 = (Gmpk85 & Nmpk85);
assign Nmpk85 = (~(vis_r0_o[14] & E5kk85));
assign Gmpk85 = (~(vis_r2_o[14] & L5kk85));
assign Slpk85 = (Umpk85 & Bnpk85);
assign Bnpk85 = (~(vis_r5_o[14] & G6kk85));
assign Umpk85 = (~(vis_r4_o[14] & N6kk85));
assign Elpk85 = (Inpk85 & Pnpk85);
assign Pnpk85 = (Wnpk85 & Dopk85);
assign Dopk85 = (~(vis_r7_o[14] & W7kk85));
assign Wnpk85 = (~(vis_r3_o[14] & D8kk85));
assign Inpk85 = (Kopk85 & Ropk85);
assign Ropk85 = (~(vis_r1_o[14] & Y8kk85));
assign Kopk85 = (~(vis_r6_o[14] & F9kk85));
assign hwdata_o[13] = (~(Sjkk85 & Yopk85));
assign Yopk85 = (Nce775 | Ubmk85);
assign Nce775 = (!Igp775);
assign Igp775 = (~(Fppk85 & Mppk85));
assign Mppk85 = (Tppk85 & Aqpk85);
assign Aqpk85 = (Hqpk85 & Oqpk85);
assign Oqpk85 = (~(vis_r11_o[13] & Eyjk85));
assign Hqpk85 = (Vqpk85 & Crpk85);
assign Crpk85 = (~(vis_r10_o[13] & Zyjk85));
assign Vqpk85 = (~(vis_r9_o[13] & Gzjk85));
assign Tppk85 = (Jrpk85 & Qrpk85);
assign Qrpk85 = (~(F3m675 & B0kk85));
assign Jrpk85 = (~(vis_r12_o[13] & I0kk85));
assign Fppk85 = (Xrpk85 & Espk85);
assign Espk85 = (Lspk85 & Sspk85);
assign Sspk85 = (~(vis_r14_o[13] & R1kk85));
assign Lspk85 = (Zspk85 & Gtpk85);
assign Gtpk85 = (~(vis_psp_o[11] & M2kk85));
assign Zspk85 = (~(vis_r8_o[13] & T2kk85));
assign Xrpk85 = (Jcy675 & Ntpk85);
assign Ntpk85 = (~(vis_msp_o[11] & H3kk85));
assign Jcy675 = (Utpk85 & Bupk85);
assign Bupk85 = (Iupk85 & Pupk85);
assign Pupk85 = (Wupk85 & Dvpk85);
assign Dvpk85 = (~(vis_r0_o[13] & E5kk85));
assign Wupk85 = (~(vis_r2_o[13] & L5kk85));
assign Iupk85 = (Kvpk85 & Rvpk85);
assign Rvpk85 = (~(vis_r5_o[13] & G6kk85));
assign Kvpk85 = (~(vis_r4_o[13] & N6kk85));
assign Utpk85 = (Yvpk85 & Fwpk85);
assign Fwpk85 = (Mwpk85 & Twpk85);
assign Twpk85 = (~(vis_r7_o[13] & W7kk85));
assign Mwpk85 = (~(vis_r3_o[13] & D8kk85));
assign Yvpk85 = (Axpk85 & Hxpk85);
assign Hxpk85 = (~(vis_r1_o[13] & Y8kk85));
assign Axpk85 = (~(vis_r6_o[13] & F9kk85));
assign Sjkk85 = (~(Ubmk85 & U7q775));
assign U7q775 = (~(Oxpk85 & Vxpk85));
assign Vxpk85 = (Cypk85 & Jypk85);
assign Jypk85 = (Qypk85 & Xypk85);
assign Xypk85 = (~(vis_r11_o[5] & Eyjk85));
assign Qypk85 = (Ezpk85 & Lzpk85);
assign Lzpk85 = (~(vis_r9_o[5] & Gzjk85));
assign Ezpk85 = (~(Asl675 & B0kk85));
assign Cypk85 = (Szpk85 & Zzpk85);
assign Zzpk85 = (~(vis_r10_o[5] & Zyjk85));
assign Szpk85 = (~(vis_psp_o[3] & M2kk85));
assign Oxpk85 = (G0qk85 & N0qk85);
assign N0qk85 = (U0qk85 & B1qk85);
assign B1qk85 = (~(vis_r12_o[5] & I0kk85));
assign U0qk85 = (I1qk85 & P1qk85);
assign P1qk85 = (~(vis_msp_o[3] & H3kk85));
assign I1qk85 = (~(vis_r14_o[5] & R1kk85));
assign G0qk85 = (E6y675 & W1qk85);
assign W1qk85 = (~(vis_r8_o[5] & T2kk85));
assign E6y675 = (D2qk85 & K2qk85);
assign K2qk85 = (R2qk85 & Y2qk85);
assign Y2qk85 = (F3qk85 & M3qk85);
assign M3qk85 = (~(vis_r0_o[5] & E5kk85));
assign F3qk85 = (~(vis_r2_o[5] & L5kk85));
assign R2qk85 = (T3qk85 & A4qk85);
assign A4qk85 = (~(vis_r5_o[5] & G6kk85));
assign T3qk85 = (~(vis_r4_o[5] & N6kk85));
assign D2qk85 = (H4qk85 & O4qk85);
assign O4qk85 = (V4qk85 & C5qk85);
assign C5qk85 = (~(vis_r7_o[5] & W7kk85));
assign V4qk85 = (~(vis_r3_o[5] & D8kk85));
assign H4qk85 = (J5qk85 & Q5qk85);
assign Q5qk85 = (~(vis_r1_o[5] & Y8kk85));
assign J5qk85 = (~(vis_r6_o[5] & F9kk85));
assign hwdata_o[12] = (~(T9kk85 & X5qk85));
assign X5qk85 = (Lie775 | Ubmk85);
assign Lie775 = (!Bgp775);
assign Bgp775 = (~(E6qk85 & L6qk85));
assign L6qk85 = (S6qk85 & Z6qk85);
assign Z6qk85 = (G7qk85 & N7qk85);
assign N7qk85 = (~(vis_r11_o[12] & Eyjk85));
assign G7qk85 = (U7qk85 & B8qk85);
assign B8qk85 = (~(vis_r9_o[12] & Gzjk85));
assign U7qk85 = (~(U1m675 & B0kk85));
assign S6qk85 = (I8qk85 & P8qk85);
assign P8qk85 = (~(vis_r10_o[12] & Zyjk85));
assign I8qk85 = (~(vis_psp_o[10] & M2kk85));
assign E6qk85 = (W8qk85 & D9qk85);
assign D9qk85 = (K9qk85 & R9qk85);
assign R9qk85 = (~(vis_r12_o[12] & I0kk85));
assign K9qk85 = (Y9qk85 & Faqk85);
assign Faqk85 = (~(vis_msp_o[10] & H3kk85));
assign Y9qk85 = (~(vis_r14_o[12] & R1kk85));
assign W8qk85 = (Qcy675 & Maqk85);
assign Maqk85 = (~(vis_r8_o[12] & T2kk85));
assign Qcy675 = (Taqk85 & Abqk85);
assign Abqk85 = (Hbqk85 & Obqk85);
assign Obqk85 = (Vbqk85 & Ccqk85);
assign Ccqk85 = (~(vis_r2_o[12] & L5kk85));
assign Vbqk85 = (~(vis_r6_o[12] & F9kk85));
assign Hbqk85 = (Jcqk85 & Qcqk85);
assign Qcqk85 = (~(vis_r5_o[12] & G6kk85));
assign Jcqk85 = (~(vis_r4_o[12] & N6kk85));
assign Taqk85 = (Xcqk85 & Edqk85);
assign Edqk85 = (Ldqk85 & Sdqk85);
assign Sdqk85 = (~(vis_r1_o[12] & Y8kk85));
assign Ldqk85 = (~(vis_r0_o[12] & E5kk85));
assign Xcqk85 = (Zdqk85 & Geqk85);
assign Geqk85 = (~(vis_r3_o[12] & D8kk85));
assign Zdqk85 = (~(vis_r7_o[12] & W7kk85));
assign T9kk85 = (~(Ubmk85 & Apq775));
assign Apq775 = (~(Neqk85 & Ueqk85));
assign Ueqk85 = (Bfqk85 & Ifqk85);
assign Ifqk85 = (Pfqk85 & Wfqk85);
assign Wfqk85 = (~(vis_r11_o[4] & Eyjk85));
assign Pfqk85 = (Dgqk85 & Kgqk85);
assign Kgqk85 = (~(vis_r9_o[4] & Gzjk85));
assign Dgqk85 = (~(Qql675 & B0kk85));
assign Bfqk85 = (Rgqk85 & Ygqk85);
assign Ygqk85 = (~(vis_r10_o[4] & Zyjk85));
assign Rgqk85 = (~(vis_psp_o[2] & M2kk85));
assign Neqk85 = (Fhqk85 & Mhqk85);
assign Mhqk85 = (Thqk85 & Aiqk85);
assign Aiqk85 = (~(vis_r12_o[4] & I0kk85));
assign Thqk85 = (Hiqk85 & Oiqk85);
assign Oiqk85 = (~(vis_msp_o[2] & H3kk85));
assign Hiqk85 = (~(vis_r14_o[4] & R1kk85));
assign Fhqk85 = (L6y675 & Viqk85);
assign Viqk85 = (~(vis_r8_o[4] & T2kk85));
assign L6y675 = (Cjqk85 & Jjqk85);
assign Jjqk85 = (Qjqk85 & Xjqk85);
assign Xjqk85 = (Ekqk85 & Lkqk85);
assign Lkqk85 = (~(vis_r0_o[4] & E5kk85));
assign Ekqk85 = (~(vis_r2_o[4] & L5kk85));
assign Qjqk85 = (Skqk85 & Zkqk85);
assign Zkqk85 = (~(vis_r5_o[4] & G6kk85));
assign Skqk85 = (~(vis_r4_o[4] & N6kk85));
assign Cjqk85 = (Glqk85 & Nlqk85);
assign Nlqk85 = (Ulqk85 & Bmqk85);
assign Bmqk85 = (~(vis_r7_o[4] & W7kk85));
assign Ulqk85 = (~(vis_r3_o[4] & D8kk85));
assign Glqk85 = (Imqk85 & Pmqk85);
assign Pmqk85 = (~(vis_r1_o[4] & Y8kk85));
assign Imqk85 = (~(vis_r6_o[4] & F9kk85));
assign hwdata_o[11] = (!Hc4775);
assign Hc4775 = (Ubmk85 ? K1d775 : Xoe775);
assign K1d775 = (!Fbp775);
assign Fbp775 = (~(Wmqk85 & Dnqk85));
assign Dnqk85 = (Knqk85 & Rnqk85);
assign Rnqk85 = (Ynqk85 & Foqk85);
assign Foqk85 = (~(vis_r11_o[3] & Eyjk85));
assign Ynqk85 = (Moqk85 & Toqk85);
assign Toqk85 = (~(vis_r9_o[3] & Gzjk85));
assign Moqk85 = (~(Gpl675 & B0kk85));
assign Knqk85 = (Apqk85 & Hpqk85);
assign Hpqk85 = (~(vis_r10_o[3] & Zyjk85));
assign Apqk85 = (~(vis_psp_o[1] & M2kk85));
assign Wmqk85 = (Opqk85 & Vpqk85);
assign Vpqk85 = (Cqqk85 & Jqqk85);
assign Jqqk85 = (~(vis_r12_o[3] & I0kk85));
assign Cqqk85 = (Qqqk85 & Xqqk85);
assign Xqqk85 = (~(vis_msp_o[1] & H3kk85));
assign Qqqk85 = (~(vis_r14_o[3] & R1kk85));
assign Opqk85 = (S6y675 & Erqk85);
assign Erqk85 = (~(vis_r8_o[3] & T2kk85));
assign S6y675 = (Lrqk85 & Srqk85);
assign Srqk85 = (Zrqk85 & Gsqk85);
assign Gsqk85 = (Nsqk85 & Usqk85);
assign Usqk85 = (~(vis_r0_o[3] & E5kk85));
assign Nsqk85 = (~(vis_r2_o[3] & L5kk85));
assign Zrqk85 = (Btqk85 & Itqk85);
assign Itqk85 = (~(vis_r5_o[3] & G6kk85));
assign Btqk85 = (~(vis_r4_o[3] & N6kk85));
assign Lrqk85 = (Ptqk85 & Wtqk85);
assign Wtqk85 = (Duqk85 & Kuqk85);
assign Kuqk85 = (~(vis_r7_o[3] & W7kk85));
assign Duqk85 = (~(vis_r3_o[3] & D8kk85));
assign Ptqk85 = (Ruqk85 & Yuqk85);
assign Yuqk85 = (~(vis_r1_o[3] & Y8kk85));
assign Ruqk85 = (~(vis_r6_o[3] & F9kk85));
assign Xoe775 = (!Wgp775);
assign Wgp775 = (~(Fvqk85 & Mvqk85));
assign Mvqk85 = (Tvqk85 & Awqk85);
assign Awqk85 = (Hwqk85 & Owqk85);
assign Owqk85 = (~(vis_r11_o[11] & Eyjk85));
assign Hwqk85 = (Vwqk85 & Cxqk85);
assign Cxqk85 = (~(vis_r10_o[11] & Zyjk85));
assign Vwqk85 = (~(vis_r9_o[11] & Gzjk85));
assign Tvqk85 = (Jxqk85 & Qxqk85);
assign Qxqk85 = (~(J0m675 & B0kk85));
assign Jxqk85 = (~(vis_r12_o[11] & I0kk85));
assign Fvqk85 = (Xxqk85 & Eyqk85);
assign Eyqk85 = (Lyqk85 & Syqk85);
assign Syqk85 = (~(vis_r14_o[11] & R1kk85));
assign Lyqk85 = (Zyqk85 & Gzqk85);
assign Gzqk85 = (~(vis_psp_o[9] & M2kk85));
assign Zyqk85 = (~(vis_r8_o[11] & T2kk85));
assign Xxqk85 = (Xcy675 & Nzqk85);
assign Nzqk85 = (~(vis_msp_o[9] & H3kk85));
assign Xcy675 = (Uzqk85 & B0rk85);
assign B0rk85 = (I0rk85 & P0rk85);
assign P0rk85 = (W0rk85 & D1rk85);
assign D1rk85 = (~(vis_r0_o[11] & E5kk85));
assign W0rk85 = (~(vis_r2_o[11] & L5kk85));
assign I0rk85 = (K1rk85 & R1rk85);
assign R1rk85 = (~(vis_r5_o[11] & G6kk85));
assign K1rk85 = (~(vis_r4_o[11] & N6kk85));
assign Uzqk85 = (Y1rk85 & F2rk85);
assign F2rk85 = (M2rk85 & T2rk85);
assign T2rk85 = (~(vis_r7_o[11] & W7kk85));
assign M2rk85 = (~(vis_r3_o[11] & D8kk85));
assign Y1rk85 = (A3rk85 & H3rk85);
assign H3rk85 = (~(vis_r1_o[11] & Y8kk85));
assign A3rk85 = (~(vis_r6_o[11] & F9kk85));
assign hwdata_o[10] = (~(J3lk85 & O3rk85));
assign O3rk85 = (Avr775 | Ubmk85);
assign Ubmk85 = (!Blkk85);
assign Avr775 = (V3rk85 & C4rk85);
assign C4rk85 = (J4rk85 & Q4rk85);
assign Q4rk85 = (X4rk85 & E5rk85);
assign E5rk85 = (~(vis_r11_o[10] & Eyjk85));
assign X4rk85 = (L5rk85 & S5rk85);
assign S5rk85 = (~(vis_r10_o[10] & Zyjk85));
assign L5rk85 = (~(vis_r9_o[10] & Gzjk85));
assign J4rk85 = (Z5rk85 & G6rk85);
assign G6rk85 = (~(Yyl675 & B0kk85));
assign Z5rk85 = (~(vis_r12_o[10] & I0kk85));
assign V3rk85 = (N6rk85 & U6rk85);
assign U6rk85 = (B7rk85 & I7rk85);
assign I7rk85 = (~(vis_r14_o[10] & R1kk85));
assign B7rk85 = (P7rk85 & W7rk85);
assign W7rk85 = (~(vis_psp_o[8] & M2kk85));
assign P7rk85 = (~(vis_r8_o[10] & T2kk85));
assign N6rk85 = (Edy675 & D8rk85);
assign D8rk85 = (~(vis_msp_o[8] & H3kk85));
assign Edy675 = (K8rk85 & R8rk85);
assign R8rk85 = (Y8rk85 & F9rk85);
assign F9rk85 = (M9rk85 & T9rk85);
assign T9rk85 = (~(vis_r0_o[10] & E5kk85));
assign M9rk85 = (~(vis_r2_o[10] & L5kk85));
assign Y8rk85 = (Aark85 & Hark85);
assign Hark85 = (~(vis_r5_o[10] & G6kk85));
assign Aark85 = (~(vis_r4_o[10] & N6kk85));
assign K8rk85 = (Oark85 & Vark85);
assign Vark85 = (Cbrk85 & Jbrk85);
assign Jbrk85 = (~(vis_r7_o[10] & W7kk85));
assign Cbrk85 = (~(vis_r3_o[10] & D8kk85));
assign Oark85 = (Qbrk85 & Xbrk85);
assign Xbrk85 = (~(vis_r1_o[10] & Y8kk85));
assign Qbrk85 = (~(vis_r6_o[10] & F9kk85));
assign J3lk85 = (Blkk85 | Neq775);
assign Neq775 = (Ecrk85 & Lcrk85);
assign Lcrk85 = (Scrk85 & Zcrk85);
assign Zcrk85 = (Gdrk85 & Ndrk85);
assign Ndrk85 = (~(Wnl675 & B0kk85));
assign Gdrk85 = (Udrk85 & Berk85);
assign Berk85 = (~(vis_psp_o[0] & M2kk85));
assign M2kk85 = (Ierk85 & Gum675);
assign Ierk85 = (Perk85 & Werk85);
assign Udrk85 = (~(vis_msp_o[0] & H3kk85));
assign H3kk85 = (Dfrk85 & Perk85);
assign Dfrk85 = (Werk85 & Kfrk85);
assign Scrk85 = (Rfrk85 & Yfrk85);
assign Yfrk85 = (~(vis_r14_o[2] & R1kk85));
assign Rfrk85 = (~(vis_r12_o[2] & I0kk85));
assign Ecrk85 = (Fgrk85 & Mgrk85);
assign Mgrk85 = (Tgrk85 & Ahrk85);
assign Ahrk85 = (~(vis_r9_o[2] & Gzjk85));
assign Tgrk85 = (Hhrk85 & Ohrk85);
assign Ohrk85 = (~(vis_r11_o[2] & Eyjk85));
assign Hhrk85 = (~(vis_r10_o[2] & Zyjk85));
assign Fgrk85 = (N7y675 & Vhrk85);
assign Vhrk85 = (~(vis_r8_o[2] & T2kk85));
assign N7y675 = (Cirk85 & Jirk85);
assign Jirk85 = (Qirk85 & Xirk85);
assign Xirk85 = (Ejrk85 & Ljrk85);
assign Ljrk85 = (~(vis_r0_o[2] & E5kk85));
assign Ejrk85 = (~(vis_r2_o[2] & L5kk85));
assign Qirk85 = (Sjrk85 & Zjrk85);
assign Zjrk85 = (~(vis_r5_o[2] & G6kk85));
assign Sjrk85 = (~(vis_r4_o[2] & N6kk85));
assign Cirk85 = (Gkrk85 & Nkrk85);
assign Nkrk85 = (Ukrk85 & Blrk85);
assign Blrk85 = (~(vis_r7_o[2] & W7kk85));
assign Ukrk85 = (~(vis_r3_o[2] & D8kk85));
assign Gkrk85 = (Ilrk85 & Plrk85);
assign Plrk85 = (~(vis_r1_o[2] & Y8kk85));
assign Ilrk85 = (~(vis_r6_o[2] & F9kk85));
assign Blkk85 = (~(Wlrk85 & Yiok85));
assign Wlrk85 = (~(Me8775 | Sunk85));
assign Me8775 = (!Oxh675);
assign hwdata_o[0] = (Oxh675 & Pgp775);
assign Pgp775 = (~(Dmrk85 & Kmrk85));
assign Kmrk85 = (Rmrk85 & Ymrk85);
assign Ymrk85 = (Fnrk85 & Mnrk85);
assign Mnrk85 = (~(vis_r10_o[0] & Zyjk85));
assign Zyjk85 = (Tnrk85 & Aork85);
assign Fnrk85 = (~(Cll675 & B0kk85));
assign B0kk85 = (Hork85 & Perk85);
assign Rmrk85 = (Oork85 & Vork85);
assign Vork85 = (~(vis_r12_o[0] & I0kk85));
assign I0kk85 = (Perk85 & Cprk85);
assign Oork85 = (~(vis_r11_o[0] & Eyjk85));
assign Eyjk85 = (Hork85 & Aork85);
assign Hork85 = (~(Bqf775 | Rgjk85));
assign Dmrk85 = (Jprk85 & Qprk85);
assign Qprk85 = (Xprk85 & Eqrk85);
assign Eqrk85 = (~(vis_r8_o[0] & T2kk85));
assign T2kk85 = (Aork85 & Cprk85);
assign Xprk85 = (~(vis_r9_o[0] & Gzjk85));
assign Gzjk85 = (Aork85 & Werk85);
assign Aork85 = (~(Yrf775 | M1i675));
assign Jprk85 = (Ldy675 & Lqrk85);
assign Lqrk85 = (~(vis_r14_o[0] & R1kk85));
assign R1kk85 = (Tnrk85 & Perk85);
assign Perk85 = (~(Yrf775 | Cnf775));
assign Tnrk85 = (~(Rgjk85 | Wyh675));
assign Ldy675 = (Sqrk85 & Zqrk85);
assign Zqrk85 = (Grrk85 & Nrrk85);
assign Nrrk85 = (Urrk85 & Bsrk85);
assign Bsrk85 = (~(vis_r0_o[0] & E5kk85));
assign E5kk85 = (Isrk85 & Cprk85);
assign Urrk85 = (~(vis_r2_o[0] & L5kk85));
assign L5kk85 = (Psrk85 & Wsrk85);
assign Psrk85 = (~(Wyh675 | M1i675));
assign Grrk85 = (Dtrk85 & Ktrk85);
assign Ktrk85 = (~(vis_r5_o[0] & G6kk85));
assign G6kk85 = (Rtrk85 & M1i675);
assign Rtrk85 = (Werk85 & Yrf775);
assign Dtrk85 = (~(vis_r4_o[0] & N6kk85));
assign N6kk85 = (Ytrk85 & M1i675);
assign Ytrk85 = (Cprk85 & Yrf775);
assign Yrf775 = (!U2i675);
assign Cprk85 = (~(Wyh675 | E0i675));
assign Sqrk85 = (Furk85 & Murk85);
assign Murk85 = (Turk85 & Avrk85);
assign Avrk85 = (~(vis_r7_o[0] & W7kk85));
assign W7kk85 = (Hvrk85 & M1i675);
assign Hvrk85 = (Wyh675 & Wsrk85);
assign Turk85 = (~(vis_r3_o[0] & D8kk85));
assign D8kk85 = (Ovrk85 & Wyh675);
assign Ovrk85 = (Wsrk85 & Cnf775);
assign Cnf775 = (!M1i675);
assign Furk85 = (Vvrk85 & Cwrk85);
assign Cwrk85 = (~(vis_r1_o[0] & Y8kk85));
assign Y8kk85 = (Isrk85 & Werk85);
assign Werk85 = (~(Bqf775 | E0i675));
assign Isrk85 = (~(M1i675 | U2i675));
assign Vvrk85 = (~(vis_r6_o[0] & F9kk85));
assign F9kk85 = (Jwrk85 & M1i675);
assign Jwrk85 = (Wsrk85 & Bqf775);
assign Bqf775 = (!Wyh675);
assign Wsrk85 = (~(Rgjk85 | U2i675));
assign Rgjk85 = (!E0i675);
assign htrans_o[1] = (Qwrk85 & Jne875);
assign Jne875 = (Prz775 | hprot_o[3]);
assign Qwrk85 = (~(Xwrk85 & Prz775));
assign Prz775 = (Exrk85 | hprot_o[0]);
assign Xwrk85 = (~(Lxrk85 & Sxrk85));
assign Sxrk85 = (Zxrk85 & Gyrk85);
assign Gyrk85 = (Fq3775 | haddr_o[28]);
assign Fq3775 = (~(Nyrk85 & haddr_o[31]));
assign Nyrk85 = (~(P8c775 | Uyrk85));
assign P8c775 = (!haddr_o[30]);
assign Zxrk85 = (~(Jlv775 | Dp3775));
assign Lxrk85 = (Yp3775 & Xl3775);
assign Yp3775 = (Bzrk85 & Qrb775);
assign Bzrk85 = (~(K61775 & Y61775));
assign K61775 = (~(B51775 & Izrk85));
assign Izrk85 = (~(Pzrk85 & O3d775));
assign hsize_o[1] = (~(Exrk85 & Wzrk85));
assign Wzrk85 = (Yiok85 | Dp3775);
assign hsize_o[0] = (D0sk85 & Sunk85);
assign D0sk85 = (Exrk85 & R61775);
assign hprot_o[3] = (~(hprot_o[2] & K0sk85));
assign K0sk85 = (~(R0sk85 & Y0sk85));
assign Y0sk85 = (~(F1sk85 & M1sk85));
assign M1sk85 = (Uyrk85 | Nx1l85[30]);
assign Uyrk85 = (!haddr_o[29]);
assign F1sk85 = (T1sk85 & A2sk85);
assign hprot_o[2] = (haddr_o[30] | haddr_o[29]);
assign haddr_o[29] = (~(H2sk85 & T1sk85));
assign T1sk85 = (Jjc775 | Gsy675);
assign Gsy675 = (Ctn775 ? O2sk85 : Cv0775);
assign O2sk85 = (V2sk85 & C3sk85);
assign C3sk85 = (J3sk85 & Q3sk85);
assign Q3sk85 = (X3sk85 & E4sk85);
assign E4sk85 = (~(Lnn775 & vis_r14_o[29]));
assign X3sk85 = (L4sk85 & S4sk85);
assign S4sk85 = (~(Gon775 & vis_psp_o[27]));
assign L4sk85 = (~(Non775 & vis_msp_o[27]));
assign J3sk85 = (Z4sk85 & G5sk85);
assign G5sk85 = (~(Ipn775 & vis_r12_o[29]));
assign Z4sk85 = (~(Ppn775 & vis_r11_o[29]));
assign V2sk85 = (N5sk85 & U5sk85);
assign U5sk85 = (B6sk85 & I6sk85);
assign I6sk85 = (~(Yqn775 & vis_r10_o[29]));
assign B6sk85 = (~(Frn775 & vis_r9_o[29]));
assign N5sk85 = (Kgy675 & P6sk85);
assign P6sk85 = (~(Trn775 & vis_r8_o[29]));
assign Kgy675 = (!E98875);
assign E98875 = (~(W6sk85 & D7sk85));
assign D7sk85 = (K7sk85 & R7sk85);
assign R7sk85 = (Y7sk85 & F8sk85);
assign F8sk85 = (~(I0c875 & vis_r0_o[29]));
assign Y7sk85 = (~(P0c875 & vis_r2_o[29]));
assign K7sk85 = (M8sk85 & T8sk85);
assign T8sk85 = (~(K1c875 & vis_r5_o[29]));
assign M8sk85 = (~(R1c875 & vis_r4_o[29]));
assign W6sk85 = (A9sk85 & H9sk85);
assign H9sk85 = (O9sk85 & V9sk85);
assign V9sk85 = (~(A3c875 & vis_r7_o[29]));
assign O9sk85 = (~(H3c875 & vis_r3_o[29]));
assign A9sk85 = (Cask85 & Jask85);
assign Jask85 = (~(C4c875 & vis_r1_o[29]));
assign Cask85 = (~(J4c875 & vis_r6_o[29]));
assign Cv0775 = (!Zpm675);
assign H2sk85 = (A2sk85 & Qask85);
assign Qask85 = (~(Nx1l85[28] & Dp3775));
assign A2sk85 = (~(Sy1l85[29] & Ms8775));
assign haddr_o[30] = (~(Xask85 & Ebsk85));
assign Ebsk85 = (~(Iq8775 & Cqy675));
assign Cqy675 = (Oln775 ? Krm675 : Lbsk85);
assign Lbsk85 = (~(Sbsk85 & Zbsk85));
assign Zbsk85 = (Gcsk85 & Ncsk85);
assign Ncsk85 = (Ucsk85 & Bdsk85);
assign Bdsk85 = (~(Lnn775 & vis_r14_o[30]));
assign Ucsk85 = (Idsk85 & Pdsk85);
assign Pdsk85 = (~(Gon775 & vis_psp_o[28]));
assign Idsk85 = (~(Non775 & vis_msp_o[28]));
assign Gcsk85 = (Wdsk85 & Desk85);
assign Desk85 = (~(Ipn775 & vis_r12_o[30]));
assign Wdsk85 = (~(Ppn775 & vis_r11_o[30]));
assign Sbsk85 = (Kesk85 & Resk85);
assign Resk85 = (Yesk85 & Ffsk85);
assign Ffsk85 = (~(Yqn775 & vis_r10_o[30]));
assign Yesk85 = (~(Frn775 & vis_r9_o[30]));
assign Kesk85 = (Wfy675 & Mfsk85);
assign Mfsk85 = (~(Trn775 & vis_r8_o[30]));
assign Wfy675 = (Tfsk85 & Agsk85);
assign Agsk85 = (Hgsk85 & Ogsk85);
assign Ogsk85 = (Vgsk85 & Chsk85);
assign Chsk85 = (~(I0c875 & vis_r0_o[30]));
assign Vgsk85 = (~(P0c875 & vis_r2_o[30]));
assign Hgsk85 = (Jhsk85 & Qhsk85);
assign Qhsk85 = (~(K1c875 & vis_r5_o[30]));
assign Jhsk85 = (~(R1c875 & vis_r4_o[30]));
assign Tfsk85 = (Xhsk85 & Eisk85);
assign Eisk85 = (Lisk85 & Sisk85);
assign Sisk85 = (~(A3c875 & vis_r7_o[30]));
assign Lisk85 = (~(H3c875 & vis_r3_o[30]));
assign Xhsk85 = (Zisk85 & Gjsk85);
assign Gjsk85 = (~(C4c875 & vis_r1_o[30]));
assign Zisk85 = (~(J4c875 & vis_r6_o[30]));
assign Xask85 = (Njsk85 & Ujsk85);
assign Ujsk85 = (~(Nx1l85[29] & Dp3775));
assign Njsk85 = (~(Sy1l85[30] & Ms8775));
assign hprot_o[0] = (~(Bksk85 & Iksk85));
assign Iksk85 = (Pksk85 & Wksk85);
assign Wksk85 = (Dlsk85 & Klsk85);
assign Dlsk85 = (Vhy775 & M2k775);
assign M2k775 = (~(Per775 & Vsg775));
assign Vhy775 = (~(Rlsk85 & Lx6775));
assign Rlsk85 = (~(Eta775 | Iso675));
assign Pksk85 = (Ylsk85 & Fmsk85);
assign Fmsk85 = (~(Mmsk85 & Oijk85));
assign Oijk85 = (Osg775 & W1p675);
assign Osg775 = (Zx6775 & X5p675);
assign Mmsk85 = (~(O6a775 | Lrh675));
assign Ylsk85 = (~(Os9775 & Tdu775));
assign Tdu775 = (X7a775 & Zry675);
assign Bksk85 = (Tmsk85 & Ansk85);
assign Ansk85 = (Hnsk85 & Jik775);
assign Hnsk85 = (R60875 & Onsk85);
assign Onsk85 = (~(Lps775 & Ub1775));
assign R60875 = (Vnsk85 & Cosk85);
assign Cosk85 = (~(Josk85 & T1s775));
assign T1s775 = (Q91775 & D1z675);
assign Josk85 = (~(F4w775 | N0p675));
assign Vnsk85 = (~(Qosk85 & Lh1775));
assign Qosk85 = (~(Te1775 | Y1z675));
assign Tmsk85 = (~(Xosk85 | X4k775));
assign X4k775 = (~(Epsk85 & Lpsk85));
assign Lpsk85 = (~(Spsk85 & A3k775));
assign Spsk85 = (~(Yyf775 | N0p675));
assign Xosk85 = (N0p675 ? Zpsk85 : Ons775);
assign Zpsk85 = (Gqsk85 & My9775);
assign Ons775 = (Vsg775 & Rto675);
assign haddr_o[7] = (~(Nqsk85 & Uqsk85));
assign Uqsk85 = (~(Nx1l85[6] & Dp3775));
assign Nqsk85 = (Brsk85 & Irsk85);
assign Irsk85 = (Jjc775 | Toy675);
assign Toy675 = (Ctn775 ? Prsk85 : E31775);
assign Prsk85 = (Wrsk85 & Dssk85);
assign Dssk85 = (Kssk85 & Rssk85);
assign Rssk85 = (Yssk85 & Ftsk85);
assign Ftsk85 = (~(Lnn775 & vis_r14_o[7]));
assign Yssk85 = (Mtsk85 & Ttsk85);
assign Ttsk85 = (~(Gon775 & vis_psp_o[5]));
assign Mtsk85 = (~(Non775 & vis_msp_o[5]));
assign Kssk85 = (Ausk85 & Husk85);
assign Husk85 = (~(Ipn775 & vis_r12_o[7]));
assign Ausk85 = (~(Ppn775 & vis_r11_o[7]));
assign Wrsk85 = (Ousk85 & Vusk85);
assign Vusk85 = (Cvsk85 & Jvsk85);
assign Jvsk85 = (~(Yqn775 & vis_r10_o[7]));
assign Cvsk85 = (~(Frn775 & vis_r9_o[7]));
assign Ousk85 = (Gey675 & Qvsk85);
assign Qvsk85 = (~(Trn775 & vis_r8_o[7]));
assign Gey675 = (!E89875);
assign E89875 = (~(Xvsk85 & Ewsk85));
assign Ewsk85 = (Lwsk85 & Swsk85);
assign Swsk85 = (Zwsk85 & Gxsk85);
assign Gxsk85 = (~(I0c875 & vis_r0_o[7]));
assign Zwsk85 = (~(P0c875 & vis_r2_o[7]));
assign Lwsk85 = (Nxsk85 & Uxsk85);
assign Uxsk85 = (~(K1c875 & vis_r5_o[7]));
assign Nxsk85 = (~(R1c875 & vis_r4_o[7]));
assign Xvsk85 = (Bysk85 & Iysk85);
assign Iysk85 = (Pysk85 & Wysk85);
assign Wysk85 = (~(A3c875 & vis_r7_o[7]));
assign Pysk85 = (~(H3c875 & vis_r3_o[7]));
assign Bysk85 = (Dzsk85 & Kzsk85);
assign Kzsk85 = (~(C4c875 & vis_r1_o[7]));
assign Dzsk85 = (~(J4c875 & vis_r6_o[7]));
assign E31775 = (!Uul675);
assign Brsk85 = (~(Sy1l85[7] & Ms8775));
assign haddr_o[6] = (~(Rzsk85 & Yzsk85));
assign Yzsk85 = (~(Nx1l85[5] & Dp3775));
assign Rzsk85 = (F0tk85 & M0tk85);
assign M0tk85 = (Jjc775 | Apy675);
assign Apy675 = (Ctn775 ? T0tk85 : Foc775);
assign T0tk85 = (A1tk85 & H1tk85);
assign H1tk85 = (O1tk85 & V1tk85);
assign V1tk85 = (C2tk85 & J2tk85);
assign J2tk85 = (~(Lnn775 & vis_r14_o[6]));
assign C2tk85 = (Q2tk85 & X2tk85);
assign X2tk85 = (~(Gon775 & vis_psp_o[4]));
assign Q2tk85 = (~(Non775 & vis_msp_o[4]));
assign O1tk85 = (E3tk85 & L3tk85);
assign L3tk85 = (~(Ipn775 & vis_r12_o[6]));
assign E3tk85 = (~(Ppn775 & vis_r11_o[6]));
assign A1tk85 = (S3tk85 & Z3tk85);
assign Z3tk85 = (G4tk85 & N4tk85);
assign N4tk85 = (~(Yqn775 & vis_r10_o[6]));
assign G4tk85 = (~(Frn775 & vis_r9_o[6]));
assign S3tk85 = (Ney675 & U4tk85);
assign U4tk85 = (~(Trn775 & vis_r8_o[6]));
assign Ney675 = (B5tk85 & I5tk85);
assign I5tk85 = (P5tk85 & W5tk85);
assign W5tk85 = (D6tk85 & K6tk85);
assign K6tk85 = (~(I0c875 & vis_r0_o[6]));
assign D6tk85 = (~(P0c875 & vis_r2_o[6]));
assign P5tk85 = (R6tk85 & Y6tk85);
assign Y6tk85 = (~(K1c875 & vis_r5_o[6]));
assign R6tk85 = (~(R1c875 & vis_r4_o[6]));
assign B5tk85 = (F7tk85 & M7tk85);
assign M7tk85 = (T7tk85 & A8tk85);
assign A8tk85 = (~(A3c875 & vis_r7_o[6]));
assign T7tk85 = (~(H3c875 & vis_r3_o[6]));
assign F7tk85 = (H8tk85 & O8tk85);
assign O8tk85 = (~(C4c875 & vis_r1_o[6]));
assign H8tk85 = (~(J4c875 & vis_r6_o[6]));
assign Foc775 = (!Ktl675);
assign F0tk85 = (~(Sy1l85[6] & Ms8775));
assign haddr_o[5] = (~(V8tk85 & C9tk85));
assign C9tk85 = (~(Nx1l85[4] & Dp3775));
assign V8tk85 = (J9tk85 & Q9tk85);
assign Q9tk85 = (Jjc775 | Hpy675);
assign Hpy675 = (Ctn775 ? X9tk85 : Duc775);
assign X9tk85 = (Eatk85 & Latk85);
assign Latk85 = (Satk85 & Zatk85);
assign Zatk85 = (Gbtk85 & Nbtk85);
assign Nbtk85 = (~(Lnn775 & vis_r14_o[5]));
assign Gbtk85 = (Ubtk85 & Bctk85);
assign Bctk85 = (~(Gon775 & vis_psp_o[3]));
assign Ubtk85 = (~(Non775 & vis_msp_o[3]));
assign Satk85 = (Ictk85 & Pctk85);
assign Pctk85 = (~(Ipn775 & vis_r12_o[5]));
assign Ictk85 = (~(Ppn775 & vis_r11_o[5]));
assign Eatk85 = (Wctk85 & Ddtk85);
assign Ddtk85 = (Kdtk85 & Rdtk85);
assign Rdtk85 = (~(Yqn775 & vis_r10_o[5]));
assign Kdtk85 = (~(Frn775 & vis_r9_o[5]));
assign Wctk85 = (Uey675 & Ydtk85);
assign Ydtk85 = (~(Trn775 & vis_r8_o[5]));
assign Uey675 = (!Lh7875);
assign Lh7875 = (~(Fetk85 & Metk85));
assign Metk85 = (Tetk85 & Aftk85);
assign Aftk85 = (Hftk85 & Oftk85);
assign Oftk85 = (~(I0c875 & vis_r0_o[5]));
assign Hftk85 = (~(P0c875 & vis_r2_o[5]));
assign Tetk85 = (Vftk85 & Cgtk85);
assign Cgtk85 = (~(K1c875 & vis_r5_o[5]));
assign Vftk85 = (~(R1c875 & vis_r4_o[5]));
assign Fetk85 = (Jgtk85 & Qgtk85);
assign Qgtk85 = (Xgtk85 & Ehtk85);
assign Ehtk85 = (~(A3c875 & vis_r7_o[5]));
assign Xgtk85 = (~(H3c875 & vis_r3_o[5]));
assign Jgtk85 = (Lhtk85 & Shtk85);
assign Shtk85 = (~(C4c875 & vis_r1_o[5]));
assign Lhtk85 = (~(J4c875 & vis_r6_o[5]));
assign Duc775 = (!Asl675);
assign J9tk85 = (~(Sy1l85[5] & Ms8775));
assign haddr_o[4] = (~(Zhtk85 & Gitk85));
assign Gitk85 = (~(Nx1l85[3] & Dp3775));
assign Zhtk85 = (Nitk85 & Uitk85);
assign Uitk85 = (Jjc775 | Opy675);
assign Opy675 = (Ctn775 ? Bjtk85 : Owc775);
assign Bjtk85 = (Ijtk85 & Pjtk85);
assign Pjtk85 = (Wjtk85 & Dktk85);
assign Dktk85 = (Kktk85 & Rktk85);
assign Rktk85 = (~(Lnn775 & vis_r14_o[4]));
assign Kktk85 = (Yktk85 & Fltk85);
assign Fltk85 = (~(Gon775 & vis_psp_o[2]));
assign Yktk85 = (~(Non775 & vis_msp_o[2]));
assign Wjtk85 = (Mltk85 & Tltk85);
assign Tltk85 = (~(Ipn775 & vis_r12_o[4]));
assign Mltk85 = (~(Ppn775 & vis_r11_o[4]));
assign Ijtk85 = (Amtk85 & Hmtk85);
assign Hmtk85 = (Omtk85 & Vmtk85);
assign Vmtk85 = (~(Yqn775 & vis_r10_o[4]));
assign Omtk85 = (~(Frn775 & vis_r9_o[4]));
assign Amtk85 = (Bfy675 & Cntk85);
assign Cntk85 = (~(Trn775 & vis_r8_o[4]));
assign Bfy675 = (!Mhb875);
assign Mhb875 = (~(Jntk85 & Qntk85));
assign Qntk85 = (Xntk85 & Eotk85);
assign Eotk85 = (Lotk85 & Sotk85);
assign Sotk85 = (~(I0c875 & vis_r0_o[4]));
assign Lotk85 = (~(P0c875 & vis_r2_o[4]));
assign Xntk85 = (Zotk85 & Gptk85);
assign Gptk85 = (~(K1c875 & vis_r5_o[4]));
assign Zotk85 = (~(R1c875 & vis_r4_o[4]));
assign Jntk85 = (Nptk85 & Uptk85);
assign Uptk85 = (Bqtk85 & Iqtk85);
assign Iqtk85 = (~(A3c875 & vis_r7_o[4]));
assign Bqtk85 = (~(H3c875 & vis_r3_o[4]));
assign Nptk85 = (Pqtk85 & Wqtk85);
assign Wqtk85 = (~(C4c875 & vis_r1_o[4]));
assign Pqtk85 = (~(J4c875 & vis_r6_o[4]));
assign Owc775 = (!Qql675);
assign Nitk85 = (~(Sy1l85[4] & Ms8775));
assign haddr_o[31] = (~(R0sk85 & Drtk85));
assign Drtk85 = (~(Nx1l85[30] & Dp3775));
assign R0sk85 = (Krtk85 & Rrtk85);
assign Rrtk85 = (Jjc775 | V2l775);
assign V2l775 = (Ctn775 ? Yrtk85 : Vlg775);
assign Yrtk85 = (Fstk85 & Mstk85);
assign Mstk85 = (Tstk85 & Attk85);
assign Attk85 = (Httk85 & Ottk85);
assign Ottk85 = (~(Lnn775 & vis_r14_o[31]));
assign Httk85 = (Vttk85 & Cutk85);
assign Cutk85 = (~(Gon775 & vis_psp_o[29]));
assign Vttk85 = (~(Non775 & vis_msp_o[29]));
assign Tstk85 = (Jutk85 & Qutk85);
assign Qutk85 = (~(Ipn775 & vis_r12_o[31]));
assign Jutk85 = (~(Ppn775 & vis_r11_o[31]));
assign Fstk85 = (Xutk85 & Evtk85);
assign Evtk85 = (Lvtk85 & Svtk85);
assign Svtk85 = (~(Yqn775 & vis_r10_o[31]));
assign Lvtk85 = (~(Frn775 & vis_r9_o[31]));
assign Xutk85 = (Pfy675 & Zvtk85);
assign Zvtk85 = (~(Trn775 & vis_r8_o[31]));
assign Pfy675 = (Gwtk85 & Nwtk85);
assign Nwtk85 = (Uwtk85 & Bxtk85);
assign Bxtk85 = (Ixtk85 & Pxtk85);
assign Pxtk85 = (~(I0c875 & vis_r0_o[31]));
assign Ixtk85 = (~(P0c875 & vis_r2_o[31]));
assign Uwtk85 = (Wxtk85 & Dytk85);
assign Dytk85 = (~(K1c875 & vis_r5_o[31]));
assign Wxtk85 = (~(R1c875 & vis_r4_o[31]));
assign Gwtk85 = (Kytk85 & Rytk85);
assign Rytk85 = (Yytk85 & Fztk85);
assign Fztk85 = (~(A3c875 & vis_r7_o[31]));
assign Yytk85 = (~(H3c875 & vis_r3_o[31]));
assign Kytk85 = (Mztk85 & Tztk85);
assign Tztk85 = (~(C4c875 & vis_r1_o[31]));
assign Mztk85 = (~(J4c875 & vis_r6_o[31]));
assign Vlg775 = (!Vsm675);
assign Krtk85 = (~(Sy1l85[31] & Ms8775));
assign haddr_o[28] = (~(A0uk85 & H0uk85));
assign H0uk85 = (~(Nx1l85[27] & Dp3775));
assign A0uk85 = (O0uk85 & V0uk85);
assign V0uk85 = (Jjc775 | Nsy675);
assign Nsy675 = (Ctn775 ? C1uk85 : V11775);
assign C1uk85 = (J1uk85 & Q1uk85);
assign Q1uk85 = (X1uk85 & E2uk85);
assign E2uk85 = (L2uk85 & S2uk85);
assign S2uk85 = (~(Lnn775 & vis_r14_o[28]));
assign L2uk85 = (Z2uk85 & G3uk85);
assign G3uk85 = (~(Gon775 & vis_psp_o[26]));
assign Z2uk85 = (~(Non775 & vis_msp_o[26]));
assign X1uk85 = (N3uk85 & U3uk85);
assign U3uk85 = (~(Ipn775 & vis_r12_o[28]));
assign N3uk85 = (~(Ppn775 & vis_r11_o[28]));
assign J1uk85 = (B4uk85 & I4uk85);
assign I4uk85 = (P4uk85 & W4uk85);
assign W4uk85 = (~(Yqn775 & vis_r10_o[28]));
assign P4uk85 = (~(Frn775 & vis_r9_o[28]));
assign B4uk85 = (Rgy675 & D5uk85);
assign D5uk85 = (~(Trn775 & vis_r8_o[28]));
assign Rgy675 = (!Y9b875);
assign Y9b875 = (~(K5uk85 & R5uk85));
assign R5uk85 = (Y5uk85 & F6uk85);
assign F6uk85 = (M6uk85 & T6uk85);
assign T6uk85 = (~(I0c875 & vis_r0_o[28]));
assign M6uk85 = (~(P0c875 & vis_r2_o[28]));
assign Y5uk85 = (A7uk85 & H7uk85);
assign H7uk85 = (~(K1c875 & vis_r5_o[28]));
assign A7uk85 = (~(R1c875 & vis_r4_o[28]));
assign K5uk85 = (O7uk85 & V7uk85);
assign V7uk85 = (C8uk85 & J8uk85);
assign J8uk85 = (~(A3c875 & vis_r7_o[28]));
assign C8uk85 = (~(H3c875 & vis_r3_o[28]));
assign O7uk85 = (Q8uk85 & X8uk85);
assign X8uk85 = (~(C4c875 & vis_r1_o[28]));
assign Q8uk85 = (~(J4c875 & vis_r6_o[28]));
assign V11775 = (!Oom675);
assign O0uk85 = (~(Sy1l85[28] & Ms8775));
assign haddr_o[27] = (~(E9uk85 & L9uk85));
assign L9uk85 = (~(Nx1l85[26] & Dp3775));
assign E9uk85 = (S9uk85 & Z9uk85);
assign Z9uk85 = (Jjc775 | Usy675);
assign Usy675 = (Ctn775 ? Gauk85 : Y9c775);
assign Gauk85 = (Nauk85 & Uauk85);
assign Uauk85 = (Bbuk85 & Ibuk85);
assign Ibuk85 = (Pbuk85 & Wbuk85);
assign Wbuk85 = (~(Lnn775 & vis_r14_o[27]));
assign Pbuk85 = (Dcuk85 & Kcuk85);
assign Kcuk85 = (~(Gon775 & vis_psp_o[25]));
assign Dcuk85 = (~(Non775 & vis_msp_o[25]));
assign Bbuk85 = (Rcuk85 & Ycuk85);
assign Ycuk85 = (~(Ipn775 & vis_r12_o[27]));
assign Rcuk85 = (~(Ppn775 & vis_r11_o[27]));
assign Nauk85 = (Fduk85 & Mduk85);
assign Mduk85 = (Tduk85 & Aeuk85);
assign Aeuk85 = (~(Yqn775 & vis_r10_o[27]));
assign Tduk85 = (~(Frn775 & vis_r9_o[27]));
assign Fduk85 = (Ygy675 & Heuk85);
assign Heuk85 = (~(Trn775 & vis_r8_o[27]));
assign Ygy675 = (!Qhd875);
assign Qhd875 = (~(Oeuk85 & Veuk85));
assign Veuk85 = (Cfuk85 & Jfuk85);
assign Jfuk85 = (Qfuk85 & Xfuk85);
assign Xfuk85 = (~(I0c875 & vis_r0_o[27]));
assign Qfuk85 = (~(P0c875 & vis_r2_o[27]));
assign Cfuk85 = (Eguk85 & Lguk85);
assign Lguk85 = (~(K1c875 & vis_r5_o[27]));
assign Eguk85 = (~(R1c875 & vis_r4_o[27]));
assign Oeuk85 = (Sguk85 & Zguk85);
assign Zguk85 = (Ghuk85 & Nhuk85);
assign Nhuk85 = (~(A3c875 & vis_r7_o[27]));
assign Ghuk85 = (~(H3c875 & vis_r3_o[27]));
assign Sguk85 = (Uhuk85 & Biuk85);
assign Biuk85 = (~(C4c875 & vis_r1_o[27]));
assign Uhuk85 = (~(J4c875 & vis_r6_o[27]));
assign Y9c775 = (!Dnm675);
assign S9uk85 = (~(Sy1l85[27] & Ms8775));
assign haddr_o[26] = (~(Iiuk85 & Piuk85));
assign Piuk85 = (~(Nx1l85[25] & Dp3775));
assign Iiuk85 = (Wiuk85 & Djuk85);
assign Djuk85 = (Jjc775 | Bty675);
assign Bty675 = (Ctn775 ? Kjuk85 : Ccc775);
assign Kjuk85 = (Rjuk85 & Yjuk85);
assign Yjuk85 = (Fkuk85 & Mkuk85);
assign Mkuk85 = (Tkuk85 & Aluk85);
assign Aluk85 = (~(Lnn775 & vis_r14_o[26]));
assign Tkuk85 = (Hluk85 & Oluk85);
assign Oluk85 = (~(Gon775 & vis_psp_o[24]));
assign Hluk85 = (~(Non775 & vis_msp_o[24]));
assign Fkuk85 = (Vluk85 & Cmuk85);
assign Cmuk85 = (~(Ipn775 & vis_r12_o[26]));
assign Vluk85 = (~(Ppn775 & vis_r11_o[26]));
assign Rjuk85 = (Jmuk85 & Qmuk85);
assign Qmuk85 = (Xmuk85 & Enuk85);
assign Enuk85 = (~(Yqn775 & vis_r10_o[26]));
assign Xmuk85 = (~(Frn775 & vis_r9_o[26]));
assign Jmuk85 = (Fhy675 & Lnuk85);
assign Lnuk85 = (~(Trn775 & vis_r8_o[26]));
assign Fhy675 = (Snuk85 & Znuk85);
assign Znuk85 = (Gouk85 & Nouk85);
assign Nouk85 = (Uouk85 & Bpuk85);
assign Bpuk85 = (~(I0c875 & vis_r0_o[26]));
assign Uouk85 = (~(P0c875 & vis_r2_o[26]));
assign Gouk85 = (Ipuk85 & Ppuk85);
assign Ppuk85 = (~(K1c875 & vis_r5_o[26]));
assign Ipuk85 = (~(R1c875 & vis_r4_o[26]));
assign Snuk85 = (Wpuk85 & Dquk85);
assign Dquk85 = (Kquk85 & Rquk85);
assign Rquk85 = (~(A3c875 & vis_r7_o[26]));
assign Kquk85 = (~(H3c875 & vis_r3_o[26]));
assign Wpuk85 = (Yquk85 & Fruk85);
assign Fruk85 = (~(C4c875 & vis_r1_o[26]));
assign Yquk85 = (~(J4c875 & vis_r6_o[26]));
assign Ccc775 = (!Slm675);
assign Wiuk85 = (~(Sy1l85[26] & Ms8775));
assign haddr_o[24] = (~(Mruk85 & Truk85));
assign Truk85 = (~(Nx1l85[23] & Dp3775));
assign Mruk85 = (Asuk85 & Hsuk85);
assign Hsuk85 = (Jjc775 | Pty675);
assign Pty675 = (Ctn775 ? Osuk85 : A20775);
assign Osuk85 = (Vsuk85 & Ctuk85);
assign Ctuk85 = (Jtuk85 & Qtuk85);
assign Qtuk85 = (Xtuk85 & Euuk85);
assign Euuk85 = (~(Lnn775 & vis_r14_o[24]));
assign Xtuk85 = (Luuk85 & Suuk85);
assign Suuk85 = (~(Gon775 & vis_psp_o[22]));
assign Luuk85 = (~(Non775 & vis_msp_o[22]));
assign Jtuk85 = (Zuuk85 & Gvuk85);
assign Gvuk85 = (~(Ipn775 & vis_r12_o[24]));
assign Zuuk85 = (~(Ppn775 & vis_r11_o[24]));
assign Vsuk85 = (Nvuk85 & Uvuk85);
assign Uvuk85 = (Bwuk85 & Iwuk85);
assign Iwuk85 = (~(Yqn775 & vis_r10_o[24]));
assign Bwuk85 = (~(Frn775 & vis_r9_o[24]));
assign Nvuk85 = (Thy675 & Pwuk85);
assign Pwuk85 = (~(Trn775 & vis_r8_o[24]));
assign Thy675 = (!C5b875);
assign C5b875 = (~(Wwuk85 & Dxuk85));
assign Dxuk85 = (Kxuk85 & Rxuk85);
assign Rxuk85 = (Yxuk85 & Fyuk85);
assign Fyuk85 = (~(I0c875 & vis_r0_o[24]));
assign Yxuk85 = (~(P0c875 & vis_r2_o[24]));
assign Kxuk85 = (Myuk85 & Tyuk85);
assign Tyuk85 = (~(K1c875 & vis_r5_o[24]));
assign Myuk85 = (~(R1c875 & vis_r4_o[24]));
assign Wwuk85 = (Azuk85 & Hzuk85);
assign Hzuk85 = (Ozuk85 & Vzuk85);
assign Vzuk85 = (~(A3c875 & vis_r7_o[24]));
assign Ozuk85 = (~(H3c875 & vis_r3_o[24]));
assign Azuk85 = (C0vk85 & J0vk85);
assign J0vk85 = (~(C4c875 & vis_r1_o[24]));
assign C0vk85 = (~(J4c875 & vis_r6_o[24]));
assign A20775 = (!Wim675);
assign Asuk85 = (~(Sy1l85[24] & Ms8775));
assign haddr_o[23] = (~(Q0vk85 & X0vk85));
assign X0vk85 = (~(Nx1l85[22] & Dp3775));
assign Q0vk85 = (E1vk85 & L1vk85);
assign L1vk85 = (Jjc775 | Wty675);
assign Wty675 = (Ctn775 ? S1vk85 : Pcf775);
assign S1vk85 = (Z1vk85 & G2vk85);
assign G2vk85 = (N2vk85 & U2vk85);
assign U2vk85 = (B3vk85 & I3vk85);
assign I3vk85 = (~(Lnn775 & vis_r14_o[23]));
assign B3vk85 = (P3vk85 & W3vk85);
assign W3vk85 = (~(Gon775 & vis_psp_o[21]));
assign P3vk85 = (~(Non775 & vis_msp_o[21]));
assign N2vk85 = (D4vk85 & K4vk85);
assign K4vk85 = (~(Ipn775 & vis_r12_o[23]));
assign D4vk85 = (~(Ppn775 & vis_r11_o[23]));
assign Z1vk85 = (R4vk85 & Y4vk85);
assign Y4vk85 = (F5vk85 & M5vk85);
assign M5vk85 = (~(Yqn775 & vis_r10_o[23]));
assign F5vk85 = (~(Frn775 & vis_r9_o[23]));
assign R4vk85 = (Aiy675 & T5vk85);
assign T5vk85 = (~(Trn775 & vis_r8_o[23]));
assign Aiy675 = (A6vk85 & H6vk85);
assign H6vk85 = (O6vk85 & V6vk85);
assign V6vk85 = (C7vk85 & J7vk85);
assign J7vk85 = (~(I0c875 & vis_r0_o[23]));
assign C7vk85 = (~(P0c875 & vis_r2_o[23]));
assign O6vk85 = (Q7vk85 & X7vk85);
assign X7vk85 = (~(K1c875 & vis_r5_o[23]));
assign Q7vk85 = (~(R1c875 & vis_r4_o[23]));
assign A6vk85 = (E8vk85 & L8vk85);
assign L8vk85 = (S8vk85 & Z8vk85);
assign Z8vk85 = (~(A3c875 & vis_r7_o[23]));
assign S8vk85 = (~(H3c875 & vis_r3_o[23]));
assign E8vk85 = (G9vk85 & N9vk85);
assign N9vk85 = (~(C4c875 & vis_r1_o[23]));
assign G9vk85 = (~(J4c875 & vis_r6_o[23]));
assign Pcf775 = (!Lhm675);
assign E1vk85 = (~(Sy1l85[23] & Ms8775));
assign haddr_o[22] = (~(U9vk85 & Bavk85));
assign Bavk85 = (~(Nx1l85[21] & Dp3775));
assign U9vk85 = (Iavk85 & Pavk85);
assign Pavk85 = (Jjc775 | Duy675);
assign Duy675 = (Ctn775 ? Wavk85 : J4d775);
assign Wavk85 = (Dbvk85 & Kbvk85);
assign Kbvk85 = (Rbvk85 & Ybvk85);
assign Ybvk85 = (Fcvk85 & Mcvk85);
assign Mcvk85 = (~(Lnn775 & vis_r14_o[22]));
assign Fcvk85 = (Tcvk85 & Advk85);
assign Advk85 = (~(Gon775 & vis_psp_o[20]));
assign Tcvk85 = (~(Non775 & vis_msp_o[20]));
assign Rbvk85 = (Hdvk85 & Odvk85);
assign Odvk85 = (~(Ipn775 & vis_r12_o[22]));
assign Hdvk85 = (~(Ppn775 & vis_r11_o[22]));
assign Dbvk85 = (Vdvk85 & Cevk85);
assign Cevk85 = (Jevk85 & Qevk85);
assign Qevk85 = (~(Yqn775 & vis_r10_o[22]));
assign Jevk85 = (~(Frn775 & vis_r9_o[22]));
assign Vdvk85 = (Hiy675 & Xevk85);
assign Xevk85 = (~(Trn775 & vis_r8_o[22]));
assign Hiy675 = (Efvk85 & Lfvk85);
assign Lfvk85 = (Sfvk85 & Zfvk85);
assign Zfvk85 = (Ggvk85 & Ngvk85);
assign Ngvk85 = (~(I0c875 & vis_r0_o[22]));
assign Ggvk85 = (~(P0c875 & vis_r2_o[22]));
assign Sfvk85 = (Ugvk85 & Bhvk85);
assign Bhvk85 = (~(K1c875 & vis_r5_o[22]));
assign Ugvk85 = (~(R1c875 & vis_r4_o[22]));
assign Efvk85 = (Ihvk85 & Phvk85);
assign Phvk85 = (Whvk85 & Divk85);
assign Divk85 = (~(A3c875 & vis_r7_o[22]));
assign Whvk85 = (~(H3c875 & vis_r3_o[22]));
assign Ihvk85 = (Kivk85 & Rivk85);
assign Rivk85 = (~(C4c875 & vis_r1_o[22]));
assign Kivk85 = (~(J4c875 & vis_r6_o[22]));
assign J4d775 = (!Agm675);
assign Iavk85 = (~(Sy1l85[22] & Ms8775));
assign haddr_o[21] = (~(Yivk85 & Fjvk85));
assign Fjvk85 = (~(Nx1l85[20] & Dp3775));
assign Yivk85 = (Mjvk85 & Tjvk85);
assign Tjvk85 = (Jjc775 | Kuy675);
assign Kuy675 = (Ctn775 ? Akvk85 : M9d775);
assign Akvk85 = (Hkvk85 & Okvk85);
assign Okvk85 = (Vkvk85 & Clvk85);
assign Clvk85 = (Jlvk85 & Qlvk85);
assign Qlvk85 = (~(Lnn775 & vis_r14_o[21]));
assign Jlvk85 = (Xlvk85 & Emvk85);
assign Emvk85 = (~(Gon775 & vis_psp_o[19]));
assign Xlvk85 = (~(Non775 & vis_msp_o[19]));
assign Vkvk85 = (Lmvk85 & Smvk85);
assign Smvk85 = (~(Ipn775 & vis_r12_o[21]));
assign Lmvk85 = (~(Ppn775 & vis_r11_o[21]));
assign Hkvk85 = (Zmvk85 & Gnvk85);
assign Gnvk85 = (Nnvk85 & Unvk85);
assign Unvk85 = (~(Yqn775 & vis_r10_o[21]));
assign Nnvk85 = (~(Frn775 & vis_r9_o[21]));
assign Zmvk85 = (Oiy675 & Bovk85);
assign Bovk85 = (~(Trn775 & vis_r8_o[21]));
assign Oiy675 = (!Ry7875);
assign Ry7875 = (~(Iovk85 & Povk85));
assign Povk85 = (Wovk85 & Dpvk85);
assign Dpvk85 = (Kpvk85 & Rpvk85);
assign Rpvk85 = (~(I0c875 & vis_r0_o[21]));
assign Kpvk85 = (~(P0c875 & vis_r2_o[21]));
assign Wovk85 = (Ypvk85 & Fqvk85);
assign Fqvk85 = (~(K1c875 & vis_r5_o[21]));
assign Ypvk85 = (~(R1c875 & vis_r4_o[21]));
assign Iovk85 = (Mqvk85 & Tqvk85);
assign Tqvk85 = (Arvk85 & Hrvk85);
assign Hrvk85 = (~(A3c875 & vis_r7_o[21]));
assign Arvk85 = (~(H3c875 & vis_r3_o[21]));
assign Mqvk85 = (Orvk85 & Vrvk85);
assign Vrvk85 = (~(C4c875 & vis_r1_o[21]));
assign Orvk85 = (~(J4c875 & vis_r6_o[21]));
assign M9d775 = (!Pem675);
assign Mjvk85 = (~(Sy1l85[21] & Ms8775));
assign haddr_o[20] = (~(Csvk85 & Jsvk85));
assign Jsvk85 = (~(Nx1l85[19] & Dp3775));
assign Csvk85 = (Qsvk85 & Xsvk85);
assign Xsvk85 = (Jjc775 | Ruy675);
assign Ruy675 = (Ctn775 ? Etvk85 : Ied775);
assign Etvk85 = (Ltvk85 & Stvk85);
assign Stvk85 = (Ztvk85 & Guvk85);
assign Guvk85 = (Nuvk85 & Uuvk85);
assign Uuvk85 = (~(Lnn775 & vis_r14_o[20]));
assign Nuvk85 = (Bvvk85 & Ivvk85);
assign Ivvk85 = (~(Gon775 & vis_psp_o[18]));
assign Bvvk85 = (~(Non775 & vis_msp_o[18]));
assign Ztvk85 = (Pvvk85 & Wvvk85);
assign Wvvk85 = (~(Ipn775 & vis_r12_o[20]));
assign Pvvk85 = (~(Ppn775 & vis_r11_o[20]));
assign Ltvk85 = (Dwvk85 & Kwvk85);
assign Kwvk85 = (Rwvk85 & Ywvk85);
assign Ywvk85 = (~(Yqn775 & vis_r10_o[20]));
assign Rwvk85 = (~(Frn775 & vis_r9_o[20]));
assign Dwvk85 = (Viy675 & Fxvk85);
assign Fxvk85 = (~(Trn775 & vis_r8_o[20]));
assign Viy675 = (!I1b875);
assign I1b875 = (~(Mxvk85 & Txvk85));
assign Txvk85 = (Ayvk85 & Hyvk85);
assign Hyvk85 = (Oyvk85 & Vyvk85);
assign Vyvk85 = (~(I0c875 & vis_r0_o[20]));
assign Oyvk85 = (~(P0c875 & vis_r2_o[20]));
assign Ayvk85 = (Czvk85 & Jzvk85);
assign Jzvk85 = (~(K1c875 & vis_r5_o[20]));
assign Czvk85 = (~(R1c875 & vis_r4_o[20]));
assign Mxvk85 = (Qzvk85 & Xzvk85);
assign Xzvk85 = (E0wk85 & L0wk85);
assign L0wk85 = (~(A3c875 & vis_r7_o[20]));
assign E0wk85 = (~(H3c875 & vis_r3_o[20]));
assign Qzvk85 = (S0wk85 & Z0wk85);
assign Z0wk85 = (~(C4c875 & vis_r1_o[20]));
assign S0wk85 = (~(J4c875 & vis_r6_o[20]));
assign Ied775 = (!Edm675);
assign Qsvk85 = (~(Sy1l85[20] & Ms8775));
assign haddr_o[1] = (~(Pzrk85 | Ckb775));
assign Ckb775 = (!O3d775);
assign O3d775 = (~(G1wk85 & N1wk85));
assign N1wk85 = (Jjc775 | Yuy675);
assign Yuy675 = (Ctn775 ? U1wk85 : Elb775);
assign U1wk85 = (B2wk85 & I2wk85);
assign I2wk85 = (P2wk85 & W2wk85);
assign W2wk85 = (D3wk85 & K3wk85);
assign K3wk85 = (~(Lnn775 & vis_r14_o[1]));
assign D3wk85 = (~(Ipn775 & vis_r12_o[1]));
assign P2wk85 = (R3wk85 & Y3wk85);
assign Y3wk85 = (~(Ppn775 & vis_r11_o[1]));
assign R3wk85 = (~(Yqn775 & vis_r10_o[1]));
assign B2wk85 = (F4wk85 & Cjy675);
assign Cjy675 = (!Bb8875);
assign Bb8875 = (~(M4wk85 & T4wk85));
assign T4wk85 = (A5wk85 & H5wk85);
assign H5wk85 = (O5wk85 & V5wk85);
assign V5wk85 = (~(I0c875 & vis_r0_o[1]));
assign O5wk85 = (~(P0c875 & vis_r2_o[1]));
assign A5wk85 = (C6wk85 & J6wk85);
assign J6wk85 = (~(K1c875 & vis_r5_o[1]));
assign C6wk85 = (~(R1c875 & vis_r4_o[1]));
assign M4wk85 = (Q6wk85 & X6wk85);
assign X6wk85 = (E7wk85 & L7wk85);
assign L7wk85 = (~(A3c875 & vis_r7_o[1]));
assign E7wk85 = (~(H3c875 & vis_r3_o[1]));
assign Q6wk85 = (S7wk85 & Z7wk85);
assign Z7wk85 = (~(C4c875 & vis_r1_o[1]));
assign S7wk85 = (~(J4c875 & vis_r6_o[1]));
assign F4wk85 = (G8wk85 & N8wk85);
assign N8wk85 = (~(Frn775 & vis_r9_o[1]));
assign G8wk85 = (~(Trn775 & vis_r8_o[1]));
assign Elb775 = (!Mml675);
assign G1wk85 = (U8wk85 & B9wk85);
assign B9wk85 = (~(Dp3775 & I9wk85));
assign I9wk85 = (~(Fj3775 ^ Ri3775));
assign Ri3775 = (!Qm2775);
assign U8wk85 = (~(Sy1l85[1] & Ms8775));
assign haddr_o[19] = (~(P9wk85 & W9wk85));
assign W9wk85 = (~(Nx1l85[18] & Dp3775));
assign P9wk85 = (Dawk85 & Kawk85);
assign Kawk85 = (Jjc775 | Fvy675);
assign Fvy675 = (Ctn775 ? Rawk85 : Ejd775);
assign Rawk85 = (Yawk85 & Fbwk85);
assign Fbwk85 = (Mbwk85 & Tbwk85);
assign Tbwk85 = (Acwk85 & Hcwk85);
assign Hcwk85 = (~(Lnn775 & vis_r14_o[19]));
assign Acwk85 = (Ocwk85 & Vcwk85);
assign Vcwk85 = (~(Gon775 & vis_psp_o[17]));
assign Ocwk85 = (~(Non775 & vis_msp_o[17]));
assign Mbwk85 = (Cdwk85 & Jdwk85);
assign Jdwk85 = (~(Ipn775 & vis_r12_o[19]));
assign Cdwk85 = (~(Ppn775 & vis_r11_o[19]));
assign Yawk85 = (Qdwk85 & Xdwk85);
assign Xdwk85 = (Eewk85 & Lewk85);
assign Lewk85 = (~(Yqn775 & vis_r10_o[19]));
assign Eewk85 = (~(Frn775 & vis_r9_o[19]));
assign Qdwk85 = (Jjy675 & Sewk85);
assign Sewk85 = (~(Trn775 & vis_r8_o[19]));
assign Jjy675 = (Zewk85 & Gfwk85);
assign Gfwk85 = (Nfwk85 & Ufwk85);
assign Ufwk85 = (Bgwk85 & Igwk85);
assign Igwk85 = (~(I0c875 & vis_r0_o[19]));
assign Bgwk85 = (~(P0c875 & vis_r2_o[19]));
assign Nfwk85 = (Pgwk85 & Wgwk85);
assign Wgwk85 = (~(K1c875 & vis_r5_o[19]));
assign Pgwk85 = (~(R1c875 & vis_r4_o[19]));
assign Zewk85 = (Dhwk85 & Khwk85);
assign Khwk85 = (Rhwk85 & Yhwk85);
assign Yhwk85 = (~(A3c875 & vis_r7_o[19]));
assign Rhwk85 = (~(H3c875 & vis_r3_o[19]));
assign Dhwk85 = (Fiwk85 & Miwk85);
assign Miwk85 = (~(C4c875 & vis_r1_o[19]));
assign Fiwk85 = (~(J4c875 & vis_r6_o[19]));
assign Ejd775 = (!Tbm675);
assign Dawk85 = (~(Sy1l85[19] & Ms8775));
assign haddr_o[18] = (~(Tiwk85 & Ajwk85));
assign Ajwk85 = (~(Nx1l85[17] & Dp3775));
assign Tiwk85 = (Hjwk85 & Ojwk85);
assign Ojwk85 = (Jjc775 | Mvy675);
assign Mvy675 = (Ctn775 ? Vjwk85 : Aod775);
assign Vjwk85 = (Ckwk85 & Jkwk85);
assign Jkwk85 = (Qkwk85 & Xkwk85);
assign Xkwk85 = (Elwk85 & Llwk85);
assign Llwk85 = (~(Lnn775 & vis_r14_o[18]));
assign Elwk85 = (Slwk85 & Zlwk85);
assign Zlwk85 = (~(Gon775 & vis_psp_o[16]));
assign Slwk85 = (~(Non775 & vis_msp_o[16]));
assign Qkwk85 = (Gmwk85 & Nmwk85);
assign Nmwk85 = (~(Ipn775 & vis_r12_o[18]));
assign Gmwk85 = (~(Ppn775 & vis_r11_o[18]));
assign Ckwk85 = (Umwk85 & Bnwk85);
assign Bnwk85 = (Inwk85 & Pnwk85);
assign Pnwk85 = (~(Yqn775 & vis_r10_o[18]));
assign Inwk85 = (~(Frn775 & vis_r9_o[18]));
assign Umwk85 = (Qjy675 & Wnwk85);
assign Wnwk85 = (~(Trn775 & vis_r8_o[18]));
assign Qjy675 = (Dowk85 & Kowk85);
assign Kowk85 = (Rowk85 & Yowk85);
assign Yowk85 = (Fpwk85 & Mpwk85);
assign Mpwk85 = (~(I0c875 & vis_r0_o[18]));
assign Fpwk85 = (~(P0c875 & vis_r2_o[18]));
assign Rowk85 = (Tpwk85 & Aqwk85);
assign Aqwk85 = (~(K1c875 & vis_r5_o[18]));
assign Tpwk85 = (~(R1c875 & vis_r4_o[18]));
assign Dowk85 = (Hqwk85 & Oqwk85);
assign Oqwk85 = (Vqwk85 & Crwk85);
assign Crwk85 = (~(A3c875 & vis_r7_o[18]));
assign Vqwk85 = (~(H3c875 & vis_r3_o[18]));
assign Hqwk85 = (Jrwk85 & Qrwk85);
assign Qrwk85 = (~(C4c875 & vis_r1_o[18]));
assign Jrwk85 = (~(J4c875 & vis_r6_o[18]));
assign Aod775 = (!Iam675);
assign Hjwk85 = (~(Sy1l85[18] & Ms8775));
assign haddr_o[17] = (~(Xrwk85 & Eswk85));
assign Eswk85 = (~(Nx1l85[16] & Dp3775));
assign Xrwk85 = (Lswk85 & Sswk85);
assign Sswk85 = (Jjc775 | Tvy675);
assign Tvy675 = (Ctn775 ? Zswk85 : Wsd775);
assign Zswk85 = (Gtwk85 & Ntwk85);
assign Ntwk85 = (Utwk85 & Buwk85);
assign Buwk85 = (Iuwk85 & Puwk85);
assign Puwk85 = (~(Lnn775 & vis_r14_o[17]));
assign Iuwk85 = (Wuwk85 & Dvwk85);
assign Dvwk85 = (~(Gon775 & vis_psp_o[15]));
assign Wuwk85 = (~(Non775 & vis_msp_o[15]));
assign Utwk85 = (Kvwk85 & Rvwk85);
assign Rvwk85 = (~(Ipn775 & vis_r12_o[17]));
assign Kvwk85 = (~(Ppn775 & vis_r11_o[17]));
assign Gtwk85 = (Yvwk85 & Fwwk85);
assign Fwwk85 = (Mwwk85 & Twwk85);
assign Twwk85 = (~(Yqn775 & vis_r10_o[17]));
assign Mwwk85 = (~(Frn775 & vis_r9_o[17]));
assign Yvwk85 = (Xjy675 & Axwk85);
assign Axwk85 = (~(Trn775 & vis_r8_o[17]));
assign Xjy675 = (!Ev7875);
assign Ev7875 = (~(Hxwk85 & Oxwk85));
assign Oxwk85 = (Vxwk85 & Cywk85);
assign Cywk85 = (Jywk85 & Qywk85);
assign Qywk85 = (~(I0c875 & vis_r0_o[17]));
assign Jywk85 = (~(P0c875 & vis_r2_o[17]));
assign Vxwk85 = (Xywk85 & Ezwk85);
assign Ezwk85 = (~(K1c875 & vis_r5_o[17]));
assign Xywk85 = (~(R1c875 & vis_r4_o[17]));
assign Hxwk85 = (Lzwk85 & Szwk85);
assign Szwk85 = (Zzwk85 & G0xk85);
assign G0xk85 = (~(A3c875 & vis_r7_o[17]));
assign Zzwk85 = (~(H3c875 & vis_r3_o[17]));
assign Lzwk85 = (N0xk85 & U0xk85);
assign U0xk85 = (~(C4c875 & vis_r1_o[17]));
assign N0xk85 = (~(J4c875 & vis_r6_o[17]));
assign Wsd775 = (!X8m675);
assign Lswk85 = (~(Sy1l85[17] & Ms8775));
assign haddr_o[15] = (~(B1xk85 & I1xk85));
assign I1xk85 = (~(Nx1l85[14] & Dp3775));
assign B1xk85 = (P1xk85 & W1xk85);
assign W1xk85 = (Jjc775 | Hwy675);
assign Hwy675 = (Ctn775 ? D2xk85 : M7f775);
assign D2xk85 = (K2xk85 & R2xk85);
assign R2xk85 = (Y2xk85 & F3xk85);
assign F3xk85 = (M3xk85 & T3xk85);
assign T3xk85 = (~(Lnn775 & vis_r14_o[15]));
assign M3xk85 = (A4xk85 & H4xk85);
assign H4xk85 = (~(Gon775 & vis_psp_o[13]));
assign A4xk85 = (~(Non775 & vis_msp_o[13]));
assign Y2xk85 = (O4xk85 & V4xk85);
assign V4xk85 = (~(Ipn775 & vis_r12_o[15]));
assign O4xk85 = (~(Ppn775 & vis_r11_o[15]));
assign K2xk85 = (C5xk85 & J5xk85);
assign J5xk85 = (Q5xk85 & X5xk85);
assign X5xk85 = (~(Yqn775 & vis_r10_o[15]));
assign Q5xk85 = (~(Frn775 & vis_r9_o[15]));
assign C5xk85 = (Lky675 & E6xk85);
assign E6xk85 = (~(Trn775 & vis_r8_o[15]));
assign Lky675 = (L6xk85 & S6xk85);
assign S6xk85 = (Z6xk85 & G7xk85);
assign G7xk85 = (N7xk85 & U7xk85);
assign U7xk85 = (~(I0c875 & vis_r0_o[15]));
assign N7xk85 = (~(P0c875 & vis_r2_o[15]));
assign Z6xk85 = (B8xk85 & I8xk85);
assign I8xk85 = (~(K1c875 & vis_r5_o[15]));
assign B8xk85 = (~(R1c875 & vis_r4_o[15]));
assign L6xk85 = (P8xk85 & W8xk85);
assign W8xk85 = (D9xk85 & K9xk85);
assign K9xk85 = (~(A3c875 & vis_r7_o[15]));
assign D9xk85 = (~(H3c875 & vis_r3_o[15]));
assign P8xk85 = (R9xk85 & Y9xk85);
assign Y9xk85 = (~(C4c875 & vis_r1_o[15]));
assign R9xk85 = (~(J4c875 & vis_r6_o[15]));
assign M7f775 = (!B6m675);
assign P1xk85 = (~(Sy1l85[15] & Ms8775));
assign haddr_o[14] = (~(Faxk85 & Maxk85));
assign Maxk85 = (~(Nx1l85[13] & Dp3775));
assign Faxk85 = (Taxk85 & Abxk85);
assign Abxk85 = (Jjc775 | Owy675);
assign Owy675 = (Ctn775 ? Hbxk85 : E4e775);
assign Hbxk85 = (Obxk85 & Vbxk85);
assign Vbxk85 = (Ccxk85 & Jcxk85);
assign Jcxk85 = (Qcxk85 & Xcxk85);
assign Xcxk85 = (~(Lnn775 & vis_r14_o[14]));
assign Qcxk85 = (Edxk85 & Ldxk85);
assign Ldxk85 = (~(Gon775 & vis_psp_o[12]));
assign Edxk85 = (~(Non775 & vis_msp_o[12]));
assign Ccxk85 = (Sdxk85 & Zdxk85);
assign Zdxk85 = (~(Ipn775 & vis_r12_o[14]));
assign Sdxk85 = (~(Ppn775 & vis_r11_o[14]));
assign Obxk85 = (Gexk85 & Nexk85);
assign Nexk85 = (Uexk85 & Bfxk85);
assign Bfxk85 = (~(Yqn775 & vis_r10_o[14]));
assign Uexk85 = (~(Frn775 & vis_r9_o[14]));
assign Gexk85 = (Sky675 & Ifxk85);
assign Ifxk85 = (~(Trn775 & vis_r8_o[14]));
assign Sky675 = (Pfxk85 & Wfxk85);
assign Wfxk85 = (Dgxk85 & Kgxk85);
assign Kgxk85 = (Rgxk85 & Ygxk85);
assign Ygxk85 = (~(I0c875 & vis_r0_o[14]));
assign Rgxk85 = (~(P0c875 & vis_r2_o[14]));
assign Dgxk85 = (Fhxk85 & Mhxk85);
assign Mhxk85 = (~(K1c875 & vis_r5_o[14]));
assign Fhxk85 = (~(R1c875 & vis_r4_o[14]));
assign Pfxk85 = (Thxk85 & Aixk85);
assign Aixk85 = (Hixk85 & Oixk85);
assign Oixk85 = (~(A3c875 & vis_r7_o[14]));
assign Hixk85 = (~(H3c875 & vis_r3_o[14]));
assign Thxk85 = (Vixk85 & Cjxk85);
assign Cjxk85 = (~(C4c875 & vis_r1_o[14]));
assign Vixk85 = (~(J4c875 & vis_r6_o[14]));
assign E4e775 = (!Q4m675);
assign Taxk85 = (~(Sy1l85[14] & Ms8775));
assign haddr_o[13] = (~(Jjxk85 & Qjxk85));
assign Qjxk85 = (~(Nx1l85[12] & Dp3775));
assign Jjxk85 = (Xjxk85 & Ekxk85);
assign Ekxk85 = (Jjc775 | Vwy675);
assign Vwy675 = (Ctn775 ? Lkxk85 : H9e775);
assign Lkxk85 = (Skxk85 & Zkxk85);
assign Zkxk85 = (Glxk85 & Nlxk85);
assign Nlxk85 = (Ulxk85 & Bmxk85);
assign Bmxk85 = (~(Lnn775 & vis_r14_o[13]));
assign Ulxk85 = (Imxk85 & Pmxk85);
assign Pmxk85 = (~(Gon775 & vis_psp_o[11]));
assign Imxk85 = (~(Non775 & vis_msp_o[11]));
assign Glxk85 = (Wmxk85 & Dnxk85);
assign Dnxk85 = (~(Ipn775 & vis_r12_o[13]));
assign Wmxk85 = (~(Ppn775 & vis_r11_o[13]));
assign Skxk85 = (Knxk85 & Rnxk85);
assign Rnxk85 = (Ynxk85 & Foxk85);
assign Foxk85 = (~(Yqn775 & vis_r10_o[13]));
assign Ynxk85 = (~(Frn775 & vis_r9_o[13]));
assign Knxk85 = (Zky675 & Moxk85);
assign Moxk85 = (~(Trn775 & vis_r8_o[13]));
assign Zky675 = (!Wq7875);
assign Wq7875 = (~(Toxk85 & Apxk85));
assign Apxk85 = (Hpxk85 & Opxk85);
assign Opxk85 = (Vpxk85 & Cqxk85);
assign Cqxk85 = (~(I0c875 & vis_r0_o[13]));
assign Vpxk85 = (~(P0c875 & vis_r2_o[13]));
assign Hpxk85 = (Jqxk85 & Qqxk85);
assign Qqxk85 = (~(K1c875 & vis_r5_o[13]));
assign Jqxk85 = (~(R1c875 & vis_r4_o[13]));
assign Toxk85 = (Xqxk85 & Erxk85);
assign Erxk85 = (Lrxk85 & Srxk85);
assign Srxk85 = (~(A3c875 & vis_r7_o[13]));
assign Lrxk85 = (~(H3c875 & vis_r3_o[13]));
assign Xqxk85 = (Zrxk85 & Gsxk85);
assign Gsxk85 = (~(C4c875 & vis_r1_o[13]));
assign Zrxk85 = (~(J4c875 & vis_r6_o[13]));
assign H9e775 = (!F3m675);
assign Xjxk85 = (~(Sy1l85[13] & Ms8775));
assign haddr_o[10] = (~(Nsxk85 & Usxk85));
assign Usxk85 = (~(Nx1l85[9] & Dp3775));
assign Dp3775 = (!R61775);
assign Nsxk85 = (Btxk85 & Itxk85);
assign Itxk85 = (Jjc775 | Qxy675);
assign Qxy675 = (Oln775 ? Nqe775 : Ptxk85);
assign Nqe775 = (!Yyl675);
assign Ptxk85 = (Wtxk85 & Duxk85);
assign Duxk85 = (Kuxk85 & Ruxk85);
assign Ruxk85 = (Yuxk85 & Fvxk85);
assign Fvxk85 = (~(Lnn775 & vis_r14_o[10]));
assign Yuxk85 = (Mvxk85 & Tvxk85);
assign Tvxk85 = (~(Gon775 & vis_psp_o[8]));
assign Gon775 = (Awxk85 & Hwxk85);
assign Awxk85 = (Owxk85 & Gum675);
assign Mvxk85 = (~(Non775 & vis_msp_o[8]));
assign Non775 = (Vwxk85 & Hwxk85);
assign Vwxk85 = (Owxk85 & Kfrk85);
assign Kfrk85 = (!Gum675);
assign Kuxk85 = (Cxxk85 & Jxxk85);
assign Jxxk85 = (~(Ipn775 & vis_r12_o[10]));
assign Cxxk85 = (~(Ppn775 & vis_r11_o[10]));
assign Wtxk85 = (Qxxk85 & Xxxk85);
assign Xxxk85 = (Eyxk85 & Lyxk85);
assign Lyxk85 = (~(Yqn775 & vis_r10_o[10]));
assign Eyxk85 = (~(Frn775 & vis_r9_o[10]));
assign Qxxk85 = (Uly675 & Syxk85);
assign Syxk85 = (~(Trn775 & vis_r8_o[10]));
assign Uly675 = (Zyxk85 & Gzxk85);
assign Gzxk85 = (Nzxk85 & Uzxk85);
assign Uzxk85 = (B0yk85 & I0yk85);
assign I0yk85 = (~(I0c875 & vis_r0_o[10]));
assign B0yk85 = (~(P0c875 & vis_r2_o[10]));
assign Nzxk85 = (P0yk85 & W0yk85);
assign W0yk85 = (~(K1c875 & vis_r5_o[10]));
assign P0yk85 = (~(R1c875 & vis_r4_o[10]));
assign Zyxk85 = (D1yk85 & K1yk85);
assign K1yk85 = (R1yk85 & Y1yk85);
assign Y1yk85 = (~(A3c875 & vis_r7_o[10]));
assign R1yk85 = (~(H3c875 & vis_r3_o[10]));
assign D1yk85 = (F2yk85 & M2yk85);
assign M2yk85 = (~(C4c875 & vis_r1_o[10]));
assign F2yk85 = (~(J4c875 & vis_r6_o[10]));
assign Btxk85 = (~(Sy1l85[10] & Ms8775));
assign haddr_o[0] = (~(Y61775 | B51775));
assign B51775 = (T2yk85 & A3yk85);
assign A3yk85 = (Jjc775 | Xxy675);
assign Xxy675 = (!Vcb775);
assign Vcb775 = (Oln775 ? Cll675 : H3yk85);
assign Oln775 = (!Ctn775);
assign Ctn775 = (O3yk85 & V3yk85);
assign V3yk85 = (C4yk85 & A7u775);
assign A7u775 = (Bbg775 | Cg8775);
assign C4yk85 = (J4yk85 & Rux775);
assign J4yk85 = (~(Q4yk85 & Hwxk85));
assign O3yk85 = (X4yk85 & E5yk85);
assign E5yk85 = (Mwo675 ? S5yk85 : L5yk85);
assign S5yk85 = (~(Sh1775 & Pw9775));
assign Sh1775 = (F6g775 & Zry675);
assign L5yk85 = (Bwg775 | Ezo675);
assign Bwg775 = (!Sa1775);
assign Sa1775 = (~(R1z675 | Rto675));
assign X4yk85 = (Z5yk85 & G6yk85);
assign G6yk85 = (~(Lfa775 & Zck775));
assign Lfa775 = (~(Ycu775 | Bvh675));
assign Z5yk85 = (~(K1z675 & N6yk85));
assign N6yk85 = (My9775 | Ub1775);
assign H3yk85 = (~(U6yk85 & B7yk85));
assign B7yk85 = (I7yk85 & P7yk85);
assign P7yk85 = (W7yk85 & D8yk85);
assign D8yk85 = (~(Lnn775 & vis_r14_o[0]));
assign Lnn775 = (Hwxk85 & Iw1l85[1]);
assign W7yk85 = (~(Ipn775 & vis_r12_o[0]));
assign Ipn775 = (Hwxk85 & K8yk85);
assign Hwxk85 = (~(Drf775 | Qnf775));
assign I7yk85 = (R8yk85 & Y8yk85);
assign Y8yk85 = (~(Ppn775 & vis_r11_o[0]));
assign Ppn775 = (Q4yk85 & F9yk85);
assign Q4yk85 = (~(Gpf775 | Vijk85));
assign R8yk85 = (~(Yqn775 & vis_r10_o[0]));
assign Yqn775 = (M9yk85 & F9yk85);
assign M9yk85 = (~(Vijk85 | Iw1l85[0]));
assign U6yk85 = (T9yk85 & Bmy675);
assign Bmy675 = (!Xjb875);
assign Xjb875 = (~(Aayk85 & Hayk85));
assign Hayk85 = (Oayk85 & Vayk85);
assign Vayk85 = (Cbyk85 & Jbyk85);
assign Jbyk85 = (~(I0c875 & vis_r0_o[0]));
assign I0c875 = (Qbyk85 & K8yk85);
assign Cbyk85 = (~(P0c875 & vis_r2_o[0]));
assign P0c875 = (Xbyk85 & Ecyk85);
assign Xbyk85 = (~(Iw1l85[0] | Iw1l85[2]));
assign Oayk85 = (Lcyk85 & Scyk85);
assign Scyk85 = (~(K1c875 & vis_r5_o[0]));
assign K1c875 = (Zcyk85 & Iw1l85[2]);
assign Zcyk85 = (Owxk85 & Drf775);
assign Lcyk85 = (~(R1c875 & vis_r4_o[0]));
assign R1c875 = (Gdyk85 & Iw1l85[2]);
assign Gdyk85 = (K8yk85 & Drf775);
assign Aayk85 = (Ndyk85 & Udyk85);
assign Udyk85 = (Beyk85 & Ieyk85);
assign Ieyk85 = (~(A3c875 & vis_r7_o[0]));
assign A3c875 = (Peyk85 & Iw1l85[2]);
assign Peyk85 = (Iw1l85[0] & Ecyk85);
assign Beyk85 = (~(H3c875 & vis_r3_o[0]));
assign H3c875 = (Weyk85 & Iw1l85[0]);
assign Weyk85 = (Ecyk85 & Qnf775);
assign Qnf775 = (!Iw1l85[2]);
assign Ndyk85 = (Dfyk85 & Kfyk85);
assign Kfyk85 = (~(C4c875 & vis_r1_o[0]));
assign C4c875 = (Qbyk85 & Owxk85);
assign Qbyk85 = (~(Iw1l85[2] | Iw1l85[3]));
assign Dfyk85 = (~(J4c875 & vis_r6_o[0]));
assign J4c875 = (Rfyk85 & Iw1l85[2]);
assign Rfyk85 = (Ecyk85 & Gpf775);
assign Ecyk85 = (~(Vijk85 | Iw1l85[3]));
assign Vijk85 = (!Iw1l85[1]);
assign T9yk85 = (Yfyk85 & Fgyk85);
assign Fgyk85 = (~(Frn775 & vis_r9_o[0]));
assign Frn775 = (F9yk85 & Owxk85);
assign Owxk85 = (~(Gpf775 | Iw1l85[1]));
assign Gpf775 = (!Iw1l85[0]);
assign Yfyk85 = (~(Trn775 & vis_r8_o[0]));
assign Trn775 = (F9yk85 & K8yk85);
assign K8yk85 = (~(Iw1l85[0] | Iw1l85[1]));
assign F9yk85 = (~(Drf775 | Iw1l85[2]));
assign Drf775 = (!Iw1l85[3]);
assign Jjc775 = (!Iq8775);
assign Iq8775 = (Mgyk85 & R61775);
assign Mgyk85 = (~(Tgyk85 & Ahyk85));
assign Ahyk85 = (Hhyk85 & Ohyk85);
assign Ohyk85 = (V1m775 | Rto675);
assign V1m775 = (!Xut775);
assign Xut775 = (R2b875 & K1z675);
assign Hhyk85 = (Vhyk85 & Ciyk85);
assign Ciyk85 = (~(Jiyk85 & Xqjk85));
assign Xqjk85 = (Rto675 & Q91775);
assign Jiyk85 = (~(Ezo675 | X5p675));
assign Vhyk85 = (Jv6875 | Ryf775);
assign Ryf775 = (!Wzr775);
assign Wzr775 = (Vxo675 & Zry675);
assign Tgyk85 = (Qiyk85 & Xiyk85);
assign Xiyk85 = (~(Yvb775 & Pw9775));
assign Qiyk85 = (Ejyk85 & Ljyk85);
assign Ljyk85 = (~(Ddt775 & U50775));
assign Ddt775 = (Ezo675 & X5p675);
assign Ejyk85 = (~(C1g775 & Mwo675));
assign C1g775 = (~(Ln9775 | K1z675));
assign T2yk85 = (~(Sy1l85[0] & Ms8775));
assign Ms8775 = (Sjyk85 & R61775);
assign R61775 = (~(Zjyk85 & Gkyk85));
assign Gkyk85 = (Nkyk85 & Ukyk85);
assign Ukyk85 = (Blyk85 & Ilyk85);
assign Ilyk85 = (~(Gqsk85 & Qza775));
assign Gqsk85 = (~(V8p675 | F3p675));
assign Blyk85 = (Plyk85 & Rny675);
assign Plyk85 = (~(O4p675 & Wlyk85));
assign Wlyk85 = (Dmyk85 | Lps775);
assign Lps775 = (D3b775 & Lh1775);
assign Dmyk85 = (Pw9775 ? Z5y775 : Yvb775);
assign Z5y775 = (Srj775 & X7a775);
assign X7a775 = (!Iso675);
assign Nkyk85 = (Kmyk85 & Rmyk85);
assign Rmyk85 = (~(Ymyk85 & Jf9775));
assign Ymyk85 = (~(K1z675 | Rto675));
assign Kmyk85 = (Fnyk85 & Mnyk85);
assign Mnyk85 = (~(Tnyk85 & Miw775));
assign Tnyk85 = (~(Te1775 | Lrh675));
assign Fnyk85 = (~(Aoyk85 & Hoyk85));
assign Aoyk85 = (Z8a775 & V0g775);
assign Zjyk85 = (Ooyk85 & Voyk85);
assign Voyk85 = (Cpyk85 & Jpyk85);
assign Jpyk85 = (~(Qpyk85 & Rvb775));
assign Qpyk85 = (~(Yaw775 | Q91775));
assign Cpyk85 = (Xpyk85 & Epsk85);
assign Epsk85 = (~(Fse875 & U50775));
assign Fse875 = (~(Ep0775 | F3p675));
assign Ep0775 = (!Vsg775);
assign Vsg775 = (Tdg775 & Cm2775);
assign Xpyk85 = (~(Eqyk85 & Lqyk85));
assign Lqyk85 = (~(Ibg775 | N0p675));
assign Eqyk85 = (~(Zry675 | Zfh775));
assign Zfh775 = (!Srj775);
assign Ooyk85 = (Sqyk85 & Jik775);
assign Jik775 = (Zqyk85 & Olg775);
assign Olg775 = (Cg8775 | K1z675);
assign Zqyk85 = (~(Zck775 & Gryk85));
assign Gryk85 = (Ps5875 | Os9775);
assign Os9775 = (Miw775 & Rto675);
assign Ps5875 = (~(Rba775 | B0z675));
assign B0z675 = (!Miw775);
assign Miw775 = (X5p675 & Pw9775);
assign Sqyk85 = (Klsk85 & Nryk85);
assign Nryk85 = (~(A3k775 & Dny675));
assign Dny675 = (~(Mwo675 | N0p675));
assign A3k775 = (Lh1775 & Cm2775);
assign Lh1775 = (~(Vya775 | V8p675));
assign Klsk85 = (Ln9775 | Y1z675);
assign Ln9775 = (!Zx6775);
assign Zx6775 = (Zry675 & Xza775);
assign Sjyk85 = (~(Uryk85 & Bsyk85));
assign Bsyk85 = (Isyk85 & Psyk85);
assign Psyk85 = (~(Fvq775 | T5a775));
assign Fvq775 = (K1z675 & Zry675);
assign Isyk85 = (Wsyk85 & Dtyk85);
assign Dtyk85 = (~(Fts775 & Psk775));
assign Fts775 = (~(Zry675 | N0p675));
assign Wsyk85 = (~(Rto675 & Ktyk85));
assign Ktyk85 = (N0p675 | Ytr775);
assign Ytr775 = (Mwo675 & Vxo675);
assign Uryk85 = (Rtyk85 & Ytyk85);
assign Ytyk85 = (Fuyk85 & Jxq775);
assign Jxq775 = (Wdl775 | Mwo675);
assign Wdl775 = (!V80875);
assign Fuyk85 = (Te1775 | Xza775);
assign Rtyk85 = (O4p675 & Muyk85);
assign Muyk85 = (Bbg775 | K1z675);
assign Y61775 = (Pzrk85 | Sunk85);
assign Sunk85 = (Yiok85 & Tuyk85);
assign Tuyk85 = (~(Avyk85 & Hvyk85));
assign Hvyk85 = (Ycu775 | W1p675);
assign Avyk85 = (~(Per775 | V80875));
assign V80875 = (Rto675 & W1p675);
assign Pzrk85 = (~(Yiok85 & Exrk85));
assign Exrk85 = (~(Ovyk85 & Vvyk85));
assign Vvyk85 = (Cl3775 & Cwyk85);
assign Cwyk85 = (~(Jwyk85 & Qwyk85));
assign Qwyk85 = (Cm2775 | Plo675);
assign Jwyk85 = (~(Jl3775 & Xwyk85));
assign Xwyk85 = (~(vis_pc_o[0] & O4y675));
assign O4y675 = (Aro675 & Exyk85);
assign Cl3775 = (Qrb775 & L40775);
assign L40775 = (!lockup_o);
assign lockup_o = (~(Lxyk85 & Sxyk85));
assign Sxyk85 = (~(Zxyk85 & Qza775));
assign Qza775 = (N0p675 & X5p675);
assign Zxyk85 = (~(M71775 | Ibg775));
assign Lxyk85 = (Gyyk85 & Nyyk85);
assign Nyyk85 = (~(Vvr775 & Uyyk85));
assign Uyyk85 = (~(Bzyk85 & Izyk85));
assign Izyk85 = (~(Pzyk85 & Wzyk85));
assign Wzyk85 = (~(Dwa775 | T17775));
assign T17775 = (!J7p675);
assign Pzyk85 = (~(Jv6875 | I6l775));
assign Jv6875 = (K7s775 | Rto675);
assign K7s775 = (!Nzy675);
assign Bzyk85 = (~(D0zk85 & Zfa775));
assign D0zk85 = (Psk775 & Y1z675);
assign Gyyk85 = (~(J7p675 & K0zk85));
assign K0zk85 = (~(Akh775 & R0zk85));
assign Akh775 = (Y0zk85 & F1zk85);
assign F1zk85 = (M1zk85 & T1zk85);
assign T1zk85 = (~(A2zk85 & H2zk85));
assign H2zk85 = (~(Yyf775 | P58775));
assign P58775 = (O2zk85 & Vbx775);
assign Vbx775 = (~(C37775 | Erj775));
assign Erj775 = (V2zk85 & C3zk85);
assign C37775 = (J3zk85 & C3zk85);
assign O2zk85 = (~(Q3zk85 | vis_primask_o));
assign Q3zk85 = (X3zk85 & E4zk85);
assign E4zk85 = (Cue875 | Ha2l85[1]);
assign Cue875 = (!Pxe875);
assign X3zk85 = (L4zk85 & Lve875);
assign Lve875 = (~(S4zk85 & Z4zk85));
assign Z4zk85 = (G5zk85 & N5zk85);
assign N5zk85 = (U5zk85 & B6zk85);
assign B6zk85 = (I6zk85 & P6zk85);
assign P6zk85 = (W6zk85 & Cb6775);
assign W6zk85 = (~(Wd7775 | Av6775));
assign I6zk85 = (~(D7zk85 | T08775));
assign U5zk85 = (K7zk85 & R7zk85);
assign R7zk85 = (~(Cq5775 | Qn8775));
assign K7zk85 = (~(Cp6775 | Xa7775));
assign G5zk85 = (Y7zk85 & F8zk85);
assign F8zk85 = (M8zk85 & T8zk85);
assign T8zk85 = (A9zk85 & V88775);
assign A9zk85 = (~(Za8775 | T9z675));
assign M8zk85 = (~(I58775 | Tm7775));
assign Y7zk85 = (H9zk85 & O9zk85);
assign O9zk85 = (~(Sj6775 | Uj7775));
assign H9zk85 = (~(P76775 | Vg7775));
assign S4zk85 = (V9zk85 & Cazk85);
assign Cazk85 = (Jazk85 & Qazk85);
assign Qazk85 = (Xazk85 & Ebzk85);
assign Ebzk85 = (Lbzk85 & B67775);
assign Lbzk85 = (~(Sbzk85 | Zbzk85));
assign Xazk85 = (~(Uti775 | Gczk85));
assign Jazk85 = (Nczk85 & Uczk85);
assign Uczk85 = (~(Jri775 | Cv7775));
assign Nczk85 = (~(Lp7775 | Qyi775));
assign V9zk85 = (Bdzk85 & Idzk85);
assign Idzk85 = (Pdzk85 & Wdzk85);
assign Wdzk85 = (~(Dd8775 | Dezk85));
assign Pdzk85 = (~(Bs6775 | Km6775));
assign Bdzk85 = (Kezk85 & Rezk85);
assign Rezk85 = (~(Yk8775 | I06775));
assign Kezk85 = (~(Rf6775 | F87775));
assign L4zk85 = (~(Yezk85 & Ffzk85));
assign Ffzk85 = (Pxe875 | G3f875);
assign G3f875 = (!Ha2l85[1]);
assign Pxe875 = (~(Mfzk85 & Tfzk85));
assign Tfzk85 = (Agzk85 & Hgzk85);
assign Hgzk85 = (Ogzk85 & Vgzk85);
assign Vgzk85 = (Chzk85 & Jhzk85);
assign Jhzk85 = (Qhzk85 & Xhzk85);
assign Xhzk85 = (Yphk85 | Gq7775);
assign Gq7775 = (!Lp7775);
assign Yphk85 = (!Mb2l85[17]);
assign Qhzk85 = (Eizk85 & Lizk85);
assign Lizk85 = (~(Ge2l85[1] & Dd8775));
assign Eizk85 = (I1jk85 | Ui8775);
assign Ui8775 = (!Dezk85);
assign I1jk85 = (!Mb2l85[35]);
assign Chzk85 = (Sizk85 & Zizk85);
assign Zizk85 = (~(Mb2l85[57] & Qyi775));
assign Sizk85 = (~(Mb2l85[49] & Jri775));
assign Ogzk85 = (Gjzk85 & Njzk85);
assign Njzk85 = (Ujzk85 & Bkzk85);
assign Bkzk85 = (Ajik85 | Xv7775);
assign Xv7775 = (!Cv7775);
assign Ajik85 = (!Mb2l85[55]);
assign Ujzk85 = (~(Mb2l85[53] & Uti775));
assign Gjzk85 = (Ikzk85 & Pkzk85);
assign Pkzk85 = (Lsik85 | Ud6775);
assign Ud6775 = (!Gczk85);
assign Lsik85 = (!Mb2l85[41]);
assign Ikzk85 = (~(Mb2l85[33] & Yk8775));
assign Agzk85 = (Wkzk85 & Dlzk85);
assign Dlzk85 = (Klzk85 & Rlzk85);
assign Rlzk85 = (Ylzk85 & Fmzk85);
assign Fmzk85 = (T3jk85 | Ey5775);
assign Ey5775 = (!Sbzk85);
assign T3jk85 = (!Mb2l85[39]);
assign Ylzk85 = (Mmzk85 & Tmzk85);
assign Tmzk85 = (~(Mb2l85[37] & I06775));
assign Mmzk85 = (L0ik85 | B67775);
assign B67775 = (!G57775);
assign L0ik85 = (!Mb2l85[31]);
assign Klzk85 = (Anzk85 & Hnzk85);
assign Hnzk85 = (X5jk85 | L56775);
assign X5jk85 = (!Mb2l85[47]);
assign Anzk85 = (~(Mb2l85[45] & P76775));
assign Wkzk85 = (Onzk85 & Vnzk85);
assign Vnzk85 = (Cozk85 & Jozk85);
assign Jozk85 = (Jshk85 | Qh7775);
assign Qh7775 = (!Vg7775);
assign Jshk85 = (!Mb2l85[23]);
assign Cozk85 = (M5hk85 | Ekj775);
assign Ekj775 = (!Sj6775);
assign M5hk85 = (!Mb2l85[15]);
assign Onzk85 = (Qozk85 & Xozk85);
assign Xozk85 = (~(Mb2l85[13] & Km6775));
assign Qozk85 = (~(Mb2l85[21] & Uj7775));
assign Mfzk85 = (Epzk85 & Lpzk85);
assign Lpzk85 = (Spzk85 & Zpzk85);
assign Zpzk85 = (Gqzk85 & Nqzk85);
assign Nqzk85 = (Uqzk85 & Brzk85);
assign Brzk85 = (Fchk85 | V88775);
assign Fchk85 = (!Mb2l85[5]);
assign Uqzk85 = (Irzk85 & Przk85);
assign Przk85 = (~(Ha2l85[1] & I58775));
assign Irzk85 = (~(Mb2l85[19] & Tm7775));
assign Gqzk85 = (Wrzk85 & Dszk85);
assign Dszk85 = (~(C92l85[1] & Rf6775));
assign Wrzk85 = (Rbhk85 | Qdi775);
assign Qdi775 = (!Za8775);
assign Rbhk85 = (!Mb2l85[3]);
assign Spzk85 = (Kszk85 & Rszk85);
assign Rszk85 = (Yszk85 & Ftzk85);
assign Ftzk85 = (~(Mb2l85[1] & T9z675));
assign Yszk85 = (~(Mb2l85[9] & Bs6775));
assign Kszk85 = (Mtzk85 & Ttzk85);
assign Ttzk85 = (I3hk85 | Xp6775);
assign Xp6775 = (!Cp6775);
assign I3hk85 = (!Mb2l85[11]);
assign Mtzk85 = (~(Mb2l85[29] & F87775));
assign Epzk85 = (Auzk85 & Huzk85);
assign Huzk85 = (Ouzk85 & Vuzk85);
assign Vuzk85 = (Cvzk85 & Jvzk85);
assign Jvzk85 = (Ayhk85 | Sb7775);
assign Sb7775 = (!Xa7775);
assign Ayhk85 = (!Mb2l85[27]);
assign Cvzk85 = (Zdjk85 | Xq5775);
assign Xq5775 = (!Cq5775);
assign Zdjk85 = (!Mb2l85[63]);
assign Ouzk85 = (Qvzk85 & Xvzk85);
assign Xvzk85 = (~(Mb2l85[61] & Qn8775));
assign Qvzk85 = (Objk85 | Wt5775);
assign Wt5775 = (!D7zk85);
assign Objk85 = (!Mb2l85[59]);
assign Auzk85 = (Ewzk85 & Lwzk85);
assign Lwzk85 = (Swzk85 & Zwzk85);
assign Zwzk85 = (Pgik85 | O18775);
assign O18775 = (!T08775);
assign Pgik85 = (!Mb2l85[51]);
assign Swzk85 = (Ssik85 | Cb6775);
assign Ssik85 = (!Mb2l85[43]);
assign Ewzk85 = (Gxzk85 & Nxzk85);
assign Nxzk85 = (~(Mb2l85[25] & Wd7775));
assign Gxzk85 = (Ybhk85 | Jcj775);
assign Ybhk85 = (!Mb2l85[7]);
assign Yezk85 = (Dye875 & N3f875);
assign N3f875 = (!Ha2l85[0]);
assign Dye875 = (~(Uxzk85 & Byzk85));
assign Byzk85 = (Iyzk85 & Pyzk85);
assign Pyzk85 = (Wyzk85 & Dzzk85);
assign Dzzk85 = (Kzzk85 & Rzzk85);
assign Rzzk85 = (Yzzk85 & F00l85);
assign F00l85 = (~(Mb2l85[16] & Lp7775));
assign Lp7775 = (~(M00l85 | T00l85));
assign Yzzk85 = (A10l85 & H10l85);
assign H10l85 = (~(Ge2l85[0] & Dd8775));
assign Dd8775 = (O10l85 & V10l85);
assign O10l85 = (C20l85 & J3zk85);
assign A10l85 = (~(Mb2l85[34] & Dezk85));
assign Dezk85 = (J20l85 & Q20l85);
assign Kzzk85 = (X20l85 & E30l85);
assign E30l85 = (~(Mb2l85[56] & Qyi775));
assign Qyi775 = (~(L30l85 | M00l85));
assign X20l85 = (~(Mb2l85[48] & Jri775));
assign Jri775 = (~(S30l85 | M00l85));
assign Wyzk85 = (Z30l85 & G40l85);
assign G40l85 = (N40l85 & U40l85);
assign U40l85 = (~(Mb2l85[54] & Cv7775));
assign Cv7775 = (B50l85 & J3zk85);
assign N40l85 = (~(Mb2l85[52] & Uti775));
assign Uti775 = (~(S30l85 | I50l85));
assign S30l85 = (!B50l85);
assign Z30l85 = (P50l85 & W50l85);
assign W50l85 = (~(Mb2l85[40] & Gczk85));
assign Gczk85 = (~(D60l85 | M00l85));
assign P50l85 = (~(Mb2l85[32] & Yk8775));
assign Yk8775 = (~(K60l85 | M00l85));
assign Iyzk85 = (R60l85 & Y60l85);
assign Y60l85 = (F70l85 & M70l85);
assign M70l85 = (T70l85 & A80l85);
assign A80l85 = (~(Mb2l85[38] & Sbzk85));
assign Sbzk85 = (J20l85 & J3zk85);
assign J20l85 = (!K60l85);
assign T70l85 = (H80l85 & O80l85);
assign O80l85 = (~(Mb2l85[36] & I06775));
assign I06775 = (~(K60l85 | I50l85));
assign K60l85 = (~(V80l85 & C90l85));
assign H80l85 = (~(Mb2l85[30] & G57775));
assign G57775 = (J90l85 & J3zk85);
assign F70l85 = (Q90l85 & X90l85);
assign X90l85 = (~(Mb2l85[46] & Zbzk85));
assign Zbzk85 = (!L56775);
assign L56775 = (D60l85 | Ea0l85);
assign Q90l85 = (~(Mb2l85[44] & P76775));
assign P76775 = (~(D60l85 | I50l85));
assign R60l85 = (La0l85 & Sa0l85);
assign Sa0l85 = (Za0l85 & Gb0l85);
assign Gb0l85 = (~(Mb2l85[22] & Vg7775));
assign Vg7775 = (J3zk85 & Nb0l85);
assign Za0l85 = (~(Mb2l85[14] & Sj6775));
assign Sj6775 = (J3zk85 & Ub0l85);
assign La0l85 = (Bc0l85 & Ic0l85);
assign Ic0l85 = (~(Mb2l85[12] & Km6775));
assign Km6775 = (~(Pc0l85 | I50l85));
assign Bc0l85 = (~(Mb2l85[20] & Uj7775));
assign Uj7775 = (~(T00l85 | I50l85));
assign T00l85 = (!Nb0l85);
assign Uxzk85 = (Wc0l85 & Dd0l85);
assign Dd0l85 = (Kd0l85 & Rd0l85);
assign Rd0l85 = (Yd0l85 & Fe0l85);
assign Fe0l85 = (Me0l85 & Te0l85);
assign Te0l85 = (S8hk85 | V88775);
assign V88775 = (Af0l85 | I50l85);
assign I50l85 = (!V2zk85);
assign S8hk85 = (!Mb2l85[4]);
assign Me0l85 = (Hf0l85 & Of0l85);
assign Of0l85 = (~(Ha2l85[0] & I58775));
assign I58775 = (Vf0l85 & Cg0l85);
assign Cg0l85 = (V10l85 & Y16775);
assign Vf0l85 = (~(Ea0l85 | Jw6775));
assign Ea0l85 = (!J3zk85);
assign Hf0l85 = (~(Mb2l85[18] & Tm7775));
assign Tm7775 = (Q20l85 & Nb0l85);
assign Nb0l85 = (Jg0l85 & vis_ipsr_o[3]);
assign Jg0l85 = (Qg0l85 & Y16775);
assign Yd0l85 = (Xg0l85 & Eh0l85);
assign Eh0l85 = (~(C92l85[0] & Rf6775));
assign Rf6775 = (Lh0l85 & V10l85);
assign Lh0l85 = (C20l85 & V2zk85);
assign Xg0l85 = (~(Mb2l85[2] & Za8775));
assign Za8775 = (Sh0l85 & Q20l85);
assign Kd0l85 = (Zh0l85 & Gi0l85);
assign Gi0l85 = (Ni0l85 & Ui0l85);
assign Ui0l85 = (~(Mb2l85[0] & T9z675));
assign T9z675 = (~(Af0l85 | M00l85));
assign Ni0l85 = (~(Mb2l85[8] & Bs6775));
assign Bs6775 = (~(Pc0l85 | M00l85));
assign M00l85 = (!Bj0l85);
assign Pc0l85 = (!Ub0l85);
assign Zh0l85 = (Ij0l85 & Pj0l85);
assign Pj0l85 = (~(Mb2l85[10] & Cp6775));
assign Cp6775 = (Ub0l85 & Q20l85);
assign Ub0l85 = (Wj0l85 & vis_ipsr_o[2]);
assign Wj0l85 = (Qg0l85 & Jw6775);
assign Ij0l85 = (~(Mb2l85[28] & F87775));
assign F87775 = (J90l85 & V2zk85);
assign Wc0l85 = (Dk0l85 & Kk0l85);
assign Kk0l85 = (Rk0l85 & Yk0l85);
assign Yk0l85 = (Fl0l85 & Ml0l85);
assign Ml0l85 = (~(Mb2l85[26] & Xa7775));
assign Xa7775 = (~(Tl0l85 | Am0l85));
assign Fl0l85 = (~(Mb2l85[62] & Cq5775));
assign Cq5775 = (Hm0l85 & J3zk85);
assign Rk0l85 = (Om0l85 & Vm0l85);
assign Vm0l85 = (~(Mb2l85[60] & Qn8775));
assign Qn8775 = (Hm0l85 & V2zk85);
assign V2zk85 = (~(Tz1775 | vis_ipsr_o[0]));
assign Om0l85 = (~(Mb2l85[58] & D7zk85));
assign D7zk85 = (Hm0l85 & Q20l85);
assign Hm0l85 = (!L30l85);
assign L30l85 = (~(C20l85 & V80l85));
assign Dk0l85 = (Cn0l85 & Jn0l85);
assign Jn0l85 = (Qn0l85 & Xn0l85);
assign Xn0l85 = (~(Mb2l85[50] & T08775));
assign T08775 = (B50l85 & Q20l85);
assign B50l85 = (Eo0l85 & V80l85);
assign Eo0l85 = (~(Jw6775 | vis_ipsr_o[2]));
assign Qn0l85 = (Kvik85 | Cb6775);
assign Cb6775 = (D60l85 | Am0l85);
assign Am0l85 = (!Q20l85);
assign Q20l85 = (~(Gw1775 | vis_ipsr_o[1]));
assign D60l85 = (~(Lo0l85 & V80l85));
assign V80l85 = (~(Ru5775 | vis_ipsr_o[4]));
assign Ru5775 = (!vis_ipsr_o[5]);
assign Lo0l85 = (~(Y16775 | vis_ipsr_o[3]));
assign Kvik85 = (!Mb2l85[42]);
assign Cn0l85 = (So0l85 & Zo0l85);
assign Zo0l85 = (~(Mb2l85[24] & Wd7775));
assign Wd7775 = (J90l85 & Bj0l85);
assign J90l85 = (!Tl0l85);
assign Tl0l85 = (~(C20l85 & Qg0l85));
assign C20l85 = (~(Y16775 | Jw6775));
assign Jw6775 = (!vis_ipsr_o[3]);
assign Y16775 = (!vis_ipsr_o[2]);
assign So0l85 = (Z8hk85 | Jcj775);
assign Jcj775 = (!Av6775);
assign Av6775 = (Sh0l85 & J3zk85);
assign J3zk85 = (~(Gw1775 | Tz1775));
assign Tz1775 = (!vis_ipsr_o[1]);
assign Gw1775 = (!vis_ipsr_o[0]);
assign Sh0l85 = (!Af0l85);
assign Af0l85 = (~(Qg0l85 & C90l85));
assign Qg0l85 = (~(Tg6775 | vis_ipsr_o[5]));
assign Tg6775 = (!vis_ipsr_o[4]);
assign Z8hk85 = (!Mb2l85[6]);
assign A2zk85 = (Z8a775 & Iah775);
assign M1zk85 = (~(Gp0l85 & Np0l85));
assign Np0l85 = (Up0l85 & Zrj775);
assign Up0l85 = (~(Ycu775 | Aay775));
assign Gp0l85 = (~(Dwa775 | Q6b775));
assign Q6b775 = (!Vvr775);
assign Dwa775 = (!Zfv775);
assign Y0zk85 = (Em3775 & Bq0l85);
assign Bq0l85 = (~(Tjh775 & Iq0l85));
assign Iq0l85 = (Pq0l85 | Wq0l85);
assign Wq0l85 = (Rpi675 ? Dr0l85 : Nc0775);
assign Dr0l85 = (~(Gwh675 | Bni675));
assign Pq0l85 = (O79775 | Cqx775);
assign Tjh775 = (Kr0l85 & Rr0l85);
assign Rr0l85 = (~(Pw9775 | Ibg775));
assign Kr0l85 = (~(I6l775 | Vya775));
assign I6l775 = (!Uag775);
assign Uag775 = (~(Xza775 | Vxo675));
assign Qrb775 = (Bav775 | Ibg775);
assign Ovyk85 = (Yr0l85 & Xl3775);
assign Xl3775 = (Fs0l85 & Ms0l85);
assign Ms0l85 = (Ts0l85 & At0l85);
assign At0l85 = (Ht0l85 & Nex775);
assign Nex775 = (Bav775 | Yyf775);
assign Yyf775 = (!T5a775);
assign T5a775 = (Q91775 & Xza775);
assign Bav775 = (~(Dba775 & Ezo675));
assign Dba775 = (X5p675 & Rto675);
assign Ht0l85 = (R0zk85 & Rny675);
assign Rny675 = (~(Vv5875 & Vvr775));
assign Vv5875 = (Ot0l85 & Ub1775);
assign Ot0l85 = (~(Del775 | U50775));
assign R0zk85 = (~(Vt0l85 & Hoyk85));
assign Hoyk85 = (~(Bbg775 | W1p675));
assign Vt0l85 = (~(R1z675 | Xuf775));
assign R1z675 = (!Rcg775);
assign Ts0l85 = (Cu0l85 & Ggh775);
assign Ggh775 = (~(Ju0l85 & Iso675));
assign Ju0l85 = (~(C8g775 | Eta775));
assign C8g775 = (!Lx6775);
assign Lx6775 = (Ezo675 & W1p675);
assign Cu0l85 = (~(Lrh675 & Qu0l85));
assign Qu0l85 = (~(Xu0l85 & Ev0l85));
assign Ev0l85 = (Lv0l85 & Sv0l85);
assign Sv0l85 = (~(Eck775 & Zv0l85));
assign Zv0l85 = (Pw9775 | Cut775);
assign Eck775 = (Z8a775 & Q91775);
assign Lv0l85 = (Gw0l85 & Att775);
assign Att775 = (~(Nw0l85 & Srj775));
assign Srj775 = (~(Eta775 | Y1z675));
assign Nw0l85 = (~(Pw9775 | U50775));
assign Gw0l85 = (~(Uw0l85 & Gvg775));
assign Uw0l85 = (~(Bvh675 | F3p675));
assign Xu0l85 = (Bx0l85 & Ix0l85);
assign Ix0l85 = (~(Gxs775 & Zfa775));
assign Bx0l85 = (Px0l85 & Wx0l85);
assign Wx0l85 = (~(Rvb775 & Dy0l85));
assign Dy0l85 = (Fjh775 | Ky0l85);
assign Ky0l85 = (~(Wnb775 | Mwo675));
assign Wnb775 = (!M7t775);
assign M7t775 = (~(Ry0l85 & Yy0l85));
assign Yy0l85 = (Fz0l85 & vis_pc_o[27]);
assign Fz0l85 = (G5i675 & Pnb775);
assign Pnb775 = (~(Bj0l85 & C3zk85));
assign C3zk85 = (V10l85 & C90l85);
assign C90l85 = (~(vis_ipsr_o[3] | vis_ipsr_o[2]));
assign V10l85 = (~(vis_ipsr_o[4] | vis_ipsr_o[5]));
assign Bj0l85 = (~(vis_ipsr_o[0] | vis_ipsr_o[1]));
assign Ry0l85 = (Mz0l85 & vis_pc_o[30]);
assign Mz0l85 = (vis_pc_o[29] & vis_pc_o[28]);
assign Rvb775 = (Z8a775 & Rto675);
assign Z8a775 = (Cm2775 & Cg8775);
assign Px0l85 = (~(Tz0l85 & Cg8775));
assign Tz0l85 = (~(A01l85 & H01l85));
assign H01l85 = (Il5875 | Xuf775);
assign Il5875 = (!D3b775);
assign D3b775 = (O01l85 & Cm2775);
assign O01l85 = (~(Ezo675 | N0p675));
assign A01l85 = (Te1775 | Y1z675);
assign Fs0l85 = (V01l85 & C11l85);
assign C11l85 = (Bqe875 & J11l85);
assign J11l85 = (~(Q11l85 & O6a775));
assign O6a775 = (X11l85 & vis_pc_o[2]);
assign X11l85 = (Doh675 & Wks775);
assign Wks775 = (!Jqh675);
assign Q11l85 = (Gxs775 & Zfa775);
assign Gxs775 = (E21l85 & My9775);
assign E21l85 = (~(Kls775 | Ezo675));
assign Kls775 = (!Rba775);
assign Rba775 = (~(L21l85 & S21l85));
assign S21l85 = (Z21l85 & G31l85);
assign G31l85 = (Ho5875 & Kc9775);
assign Kc9775 = (Bx8775 | Amf775);
assign Bx8775 = (!N1j675);
assign Ho5875 = (~(J0j675 & C27875));
assign C27875 = (Y3b775 | Fzi675);
assign Z21l85 = (Ncz775 & Km5875);
assign Km5875 = (~(Fzi675 & Y3b775));
assign Y3b775 = (N31l85 | Byi675);
assign Ncz775 = (~(Byi675 & N31l85));
assign N31l85 = (!M86875);
assign M86875 = (F4b775 & N1p775);
assign L21l85 = (U31l85 & B41l85);
assign B41l85 = (~(R2j675 & I41l85));
assign I41l85 = (V3j675 | N1j675);
assign U31l85 = (Gv9775 & C5x775);
assign C5x775 = (N1p775 | F4b775);
assign F4b775 = (!Pl5875);
assign Pl5875 = (T4b775 | A5j675);
assign N1p775 = (!Xwi675);
assign Gv9775 = (~(A5j675 & T4b775));
assign T4b775 = (~(P41l85 & Amf775));
assign Amf775 = (!V3j675);
assign P41l85 = (~(N1j675 | R2j675));
assign Bqe875 = (!Fyg775);
assign Fyg775 = (Rcg775 & My9775);
assign Rcg775 = (~(Xza775 | N0p675));
assign V01l85 = (W41l85 & D51l85);
assign D51l85 = (~(Nzy675 & Rfr775));
assign W41l85 = (N0p675 ? R51l85 : K51l85);
assign R51l85 = (M71775 | Ibg775);
assign K51l85 = (Y51l85 & F61l85);
assign F61l85 = (~(Yvb775 & Ub1775));
assign Y51l85 = (M61l85 & T61l85);
assign T61l85 = (~(A71l85 & Iso675));
assign A71l85 = (~(Za1775 | Eta775));
assign M61l85 = (~(Per775 & My9775));
assign Per775 = (Q91775 & U50775);
assign Yr0l85 = (Em3775 & H71l85);
assign H71l85 = (~(O71l85 & Fj3775));
assign Fj3775 = (!vis_pc_o[0]);
assign O71l85 = (~(Jl3775 & Qm2775));
assign Qm2775 = (~(Spo675 & Exyk85));
assign Exyk85 = (F80775 | Fg5875);
assign F80775 = (~(Vtt775 | V71l85));
assign V71l85 = (Frg775 & K1z675);
assign Frg775 = (~(Q91775 | Bvh675));
assign Vtt775 = (Jf9775 & Mwo675);
assign Jl3775 = (H90775 | Fg5875);
assign Fg5875 = (C81l85 & J81l85);
assign J81l85 = (Q81l85 & X81l85);
assign X81l85 = (E91l85 & L91l85);
assign L91l85 = (~(S91l85 & Z91l85));
assign Z91l85 = (~(Ycu775 | Q91775));
assign Ycu775 = (!Oay775);
assign Oay775 = (~(Xza775 | Rto675));
assign S91l85 = (~(Veg775 | E5z675));
assign Veg775 = (!M4w775);
assign M4w775 = (~(W1p675 | O4p675));
assign E91l85 = (Ga1l85 & Ncl775);
assign Ncl775 = (Mbw775 | Nvg775);
assign Nvg775 = (!M6g775);
assign M6g775 = (~(Q91775 | O4p675));
assign Mbw775 = (!T2r775);
assign T2r775 = (W1p675 & Xza775);
assign Ga1l85 = (~(Na1l85 & Ua1l85));
assign Ua1l85 = (Kny675 & Xza775);
assign Na1l85 = (~(Bbg775 | Sn9775));
assign Sn9775 = (E5z675 | Rto675);
assign Q81l85 = (Bb1l85 & Ib1l85);
assign Ib1l85 = (~(Pb1l85 & Lsw775));
assign Lsw775 = (~(Vya775 | Y1z675));
assign Vya775 = (!Eew775);
assign Pb1l85 = (Wb1l85 & Te1775);
assign Te1775 = (!Zck775);
assign Zck775 = (W1p675 & Zry675);
assign Wb1l85 = (Zfa775 | Iah775);
assign Iah775 = (K1z675 & U50775);
assign Zfa775 = (K1z675 & Pw9775);
assign Bb1l85 = (~(Dc1l85 & Xxq775));
assign Xxq775 = (W1p675 & D1z675);
assign D1z675 = (!O4p675);
assign Dc1l85 = (~(Y1z675 | X5p675));
assign C81l85 = (Kc1l85 & Rc1l85);
assign Rc1l85 = (Yc1l85 & Fd1l85);
assign Fd1l85 = (~(Md1l85 & Psk775));
assign Psk775 = (~(W1p675 | X5p675));
assign Md1l85 = (V0g775 & Vvr775);
assign Vvr775 = (~(Zry675 | Bvh675));
assign V0g775 = (~(Vxo675 | F3p675));
assign Yc1l85 = (~(J7p675 & Td1l85));
assign Td1l85 = (~(Em3775 & Ae1l85));
assign Ae1l85 = (~(He1l85 & Gvg775));
assign Gvg775 = (Vxo675 & U50775);
assign He1l85 = (~(Xuf775 | Bbg775));
assign Kc1l85 = (Oe1l85 & Ve1l85);
assign Ve1l85 = (~(Gwf775 & Cf1l85));
assign Cf1l85 = (~(Jf1l85 & Qf1l85));
assign Qf1l85 = (~(T0m775 | O4p675));
assign Jf1l85 = (~(Fjh775 | Nzy675));
assign Nzy675 = (Mwo675 & U50775);
assign Fjh775 = (Vxo675 & Pw9775);
assign Pw9775 = (!N0p675);
assign Gwf775 = (Bvh675 & M71775);
assign Oe1l85 = (~(N0p675 & Xf1l85));
assign Xf1l85 = (~(Eg1l85 & Lg1l85));
assign Lg1l85 = (Sg1l85 & Zg1l85);
assign Zg1l85 = (~(Unv775 | Yvb775));
assign Yvb775 = (F6g775 & R2b875);
assign F6g775 = (W1p675 & K1z675);
assign Unv775 = (My9775 & F3p675);
assign Sg1l85 = (Gh1l85 & Nh1l85);
assign Nh1l85 = (~(J7p675 & Uh1l85));
assign Uh1l85 = (~(Bi1l85 & Ii1l85));
assign Ii1l85 = (~(Mjh775 & Eew775));
assign Mjh775 = (~(Bbg775 | Rpi675));
assign Bbg775 = (!R2b875);
assign R2b875 = (~(Zry675 | Q91775));
assign Bi1l85 = (~(Pi1l85 & Y1z675));
assign Pi1l85 = (~(Wi1l85 & Dj1l85));
assign Dj1l85 = (~(Kj1l85 & Zfv775));
assign Zfv775 = (~(Lrh675 | Rpi675));
assign Kj1l85 = (~(Zry675 | Aay775));
assign Aay775 = (Ilk775 & Rj1l85);
assign Rj1l85 = (Ty2775 | Iw2775);
assign Iw2775 = (!Vci675);
assign Ty2775 = (!Cei675);
assign Ilk775 = (Jfi675 & Iq1775);
assign Iq1775 = (!Qgi675);
assign Wi1l85 = (~(Eew775 & Yj1l85));
assign Yj1l85 = (~(Fk1l85 & Dhw775));
assign Dhw775 = (Ryt775 & Mk1l85);
assign Mk1l85 = (Rpi675 | Zqi675);
assign Ryt775 = (!Cqx775);
assign Cqx775 = (Bni675 & Hk3775);
assign Hk3775 = (!Rpi675);
assign Fk1l85 = (Tk1l85 & Jqx775);
assign Jqx775 = (!O79775);
assign O79775 = (E2u775 & Nc0775);
assign E2u775 = (!Gwh675);
assign Tk1l85 = (~(Rpi675 & Hay775));
assign Hay775 = (~(Nc0775 | Bni675));
assign Nc0775 = (!Zqi675);
assign Eew775 = (~(Lrh675 | X5p675));
assign Gh1l85 = (Za1775 | Eta775);
assign Eta775 = (!Rfr775);
assign Rfr775 = (~(Cg8775 | Xza775));
assign Xza775 = (!F3p675);
assign Za1775 = (!Gtb775);
assign Gtb775 = (Zry675 & U50775);
assign Zry675 = (!Ezo675);
assign Eg1l85 = (~(Al1l85 | Hl1l85));
assign Hl1l85 = (V8p675 ? My9775 : Ol1l85);
assign My9775 = (X5p675 & Y1z675);
assign Ol1l85 = (~(Xuf775 | K1z675));
assign Al1l85 = (~(Vl1l85 & Cm1l85));
assign Cm1l85 = (Yaw775 | U3g775);
assign U3g775 = (!Cut775);
assign Cut775 = (W1p675 & Y1z675);
assign Yaw775 = (!Wc1775);
assign Wc1775 = (E5z675 & M71775);
assign M71775 = (!V8p675);
assign E5z675 = (!Lrh675);
assign Vl1l85 = (F4w775 | Q91775);
assign F4w775 = (!Tdg775);
assign Tdg775 = (~(K1z675 | Lrh675));
assign H90775 = (Rux775 & Jm1l85);
assign Jm1l85 = (~(Nsx775 & W1p675));
assign Nsx775 = (~(Oya775 | Mwo675));
assign Oya775 = (!Jf9775);
assign Jf9775 = (N0p675 & Cm2775);
assign Cm2775 = (!Bvh675);
assign Rux775 = (!Z8v775);
assign Z8v775 = (Zrj775 & X5p675);
assign Zrj775 = (N0p675 & Q91775);
assign Em3775 = (Lbz775 & Qm1l85);
assign Qm1l85 = (~(Pzr775 & Jlv775));
assign Pzr775 = (~(Y1z675 | Q91775));
assign Lbz775 = (Xuf775 | Kp3775);
assign Kp3775 = (!Jlv775);
assign Jlv775 = (V8p675 & Cg8775);
assign Cg8775 = (!X5p675);
assign Xuf775 = (!Ub1775);
assign Ub1775 = (O4p675 & Y1z675);
assign Y1z675 = (!Rto675);
assign Yiok85 = (Xm1l85 & En1l85);
assign En1l85 = (Ln1l85 & Duq775);
assign Duq775 = (!Fku775);
assign Fku775 = (Q91775 & K1z675);
assign K1z675 = (!Vxo675);
assign Ln1l85 = (~(Sn1l85 & F3p675));
assign Sn1l85 = (Mwo675 & Kny675);
assign Kny675 = (Vxo675 & W1p675);
assign Xm1l85 = (Zn1l85 & Go1l85);
assign Go1l85 = (Ibg775 | Del775);
assign Del775 = (!T0m775);
assign T0m775 = (F3p675 & Q91775);
assign Q91775 = (!Mwo675);
assign Ibg775 = (!Rtr775);
assign Rtr775 = (O4p675 & U50775);
assign U50775 = (!W1p675);
assign Zn1l85 = (Ezo675 | Bvh675);

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ih3l85 <= 1'b0;
  else
    Ih3l85 <= D2y675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yi3l85 <= 1'b1;
  else
    Yi3l85 <= G0y675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gk3l85 <= 1'b1;
  else
    Gk3l85 <= Elx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vl3l85 <= 1'b1;
  else
    Vl3l85 <= Y1s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fn3l85 <= 1'b1;
  else
    Fn3l85 <= H3s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Oo3l85 <= 1'b1;
  else
    Oo3l85 <= R1s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yp3l85 <= 1'b0;
  else
    Yp3l85 <= Xyx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hr3l85 <= 1'b1;
  else
    Hr3l85 <= Oev675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qs3l85 <= 1'b1;
  else
    Qs3l85 <= Hev675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fu3l85 <= 1'b0;
  else
    Fu3l85 <= Cyq675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xv3l85 <= 1'b0;
  else
    Xv3l85 <= T2s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kx3l85 <= 1'b0;
  else
    Kx3l85 <= K1s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vy3l85 <= 1'b0;
  else
    Vy3l85 <= D1s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I04l85 <= 1'b1;
  else
    I04l85 <= W0s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    W14l85 <= 1'b1;
  else
    W14l85 <= N6s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    L34l85 <= 1'b0;
  else
    L34l85 <= Ggw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Z44l85 <= 1'b1;
  else
    Z44l85 <= Rqv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    O64l85 <= 1'b1;
  else
    O64l85 <= Oxx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    D84l85 <= 1'b0;
  else
    D84l85 <= Szq675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    V94l85 <= 1'b1;
  else
    V94l85 <= Dqv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jb4l85 <= 1'b1;
  else
    Jb4l85 <= Axx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xc4l85 <= 1'b0;
  else
    Xc4l85 <= W9q675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pe4l85 <= 1'b1;
  else
    Pe4l85 <= Ntx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dg4l85 <= 1'b1;
  else
    Dg4l85 <= Iux675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rh4l85 <= 1'b1;
  else
    Rh4l85 <= Lzx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fj4l85 <= 1'b1;
  else
    Fj4l85 <= Wpv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tk4l85 <= 1'b1;
  else
    Tk4l85 <= Ezx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hm4l85 <= 1'b0;
  else
    Hm4l85 <= Aqq675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zn4l85 <= 1'b1;
  else
    Zn4l85 <= Ssx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kp4l85 <= 1'b1;
  else
    Kp4l85 <= Hlv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yq4l85 <= 1'b0;
  else
    Yq4l85 <= J9u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Os4l85 <= 1'b1;
  else
    Os4l85 <= Sbt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Du4l85 <= 1'b1;
  else
    Du4l85 <= Uct675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sv4l85 <= 1'b0;
  else
    Sv4l85 <= G8q675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kx4l85 <= 1'b1;
  else
    Kx4l85 <= P0s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wy4l85 <= 1'b0;
  else
    Wy4l85 <= I0s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    J05l85 <= 1'b0;
  else
    J05l85 <= B0s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    W15l85 <= 1'b1;
  else
    W15l85 <= Uzr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    K35l85 <= 1'b1;
  else
    K35l85 <= Znv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Z45l85 <= 1'b1;
  else
    Z45l85 <= Lnv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    N65l85 <= 1'b1;
  else
    N65l85 <= Env675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    B85l85 <= 1'b1;
  else
    B85l85 <= Ebt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Q95l85 <= 1'b1;
  else
    Q95l85 <= Yvx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fb5l85 <= 1'b1;
  else
    Fb5l85 <= Kvx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tc5l85 <= 1'b1;
  else
    Tc5l85 <= Dvx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    He5l85 <= 1'b1;
  else
    He5l85 <= A9t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wf5l85 <= 1'b1;
  else
    Wf5l85 <= V3s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lh5l85 <= 1'b0;
  else
    Lh5l85 <= M3y675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bj5l85 <= 1'b1;
  else
    Bj5l85 <= Fsu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qk5l85 <= 1'b1;
  else
    Qk5l85 <= Juu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fm5l85 <= 1'b1;
  else
    Fm5l85 <= Xuu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Un5l85 <= 1'b1;
  else
    Un5l85 <= Zvu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jp5l85 <= 1'b0;
  else
    Jp5l85 <= Koq675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Br5l85 <= 1'b1;
  else
    Br5l85 <= Lsx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ps5l85 <= 1'b1;
  else
    Ps5l85 <= G2w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Du5l85 <= 1'b0;
  else
    Du5l85 <= Alv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ov5l85 <= 1'b1;
  else
    Ov5l85 <= Dms675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cx5l85 <= 1'b1;
  else
    Cx5l85 <= Hos675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qy5l85 <= 1'b1;
  else
    Qy5l85 <= Vos675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    E06l85 <= 1'b1;
  else
    E06l85 <= Xps675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    S16l85 <= 1'b0;
  else
    S16l85 <= U1q675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    K36l85 <= 1'b0;
  else
    K36l85 <= Vdw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    V46l85 <= 1'b1;
  else
    V46l85 <= Nzr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    G66l85 <= 1'b1;
  else
    G66l85 <= K2y675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    V76l85 <= 1'b0;
  else
    V76l85 <= Gzr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I96l85 <= 1'b0;
  else
    I96l85 <= Zyr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Va6l85 <= 1'b1;
  else
    Va6l85 <= Syr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fc6l85 <= 1'b0;
  else
    Fc6l85 <= Lyr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vd6l85 <= 1'b0;
  else
    Vd6l85 <= U9w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hf6l85 <= 1'b1;
  else
    Hf6l85 <= R2y675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wg6l85 <= 1'b1;
  else
    Wg6l85 <= Fpx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Li6l85 <= 1'b1;
  else
    Li6l85 <= Yox675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ak6l85 <= 1'b0;
  else
    Ak6l85 <= Rox675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ml6l85 <= 1'b1;
  else
    Ml6l85 <= Zzx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bn6l85 <= 1'b1;
  else
    Bn6l85 <= Eyr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Po6l85 <= 1'b1;
  else
    Po6l85 <= Meu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dq6l85 <= 1'b1;
  else
    Dq6l85 <= Qgu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rr6l85 <= 1'b1;
  else
    Rr6l85 <= Ehu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ft6l85 <= 1'b1;
  else
    Ft6l85 <= Giu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tu6l85 <= 1'b0;
  else
    Tu6l85 <= Yhq675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lw6l85 <= 1'b0;
  else
    Lw6l85 <= Jyx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ux6l85 <= 1'b1;
  else
    Ux6l85 <= Snv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jz6l85 <= 1'b1;
  else
    Jz6l85 <= Kqv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Y07l85 <= 1'b1;
  else
    Y07l85 <= Rvx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    N27l85 <= 1'b1;
  else
    N27l85 <= Vxx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    C47l85 <= 1'b0;
  else
    C47l85 <= Wuq675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    U57l85 <= 1'b0;
  else
    U57l85 <= Fcw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    F77l85 <= 1'b1;
  else
    F77l85 <= Niu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    T87l85 <= 1'b0;
  else
    T87l85 <= I1y675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ja7l85 <= 1'b1;
  else
    Ja7l85 <= K8s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yb7l85 <= 1'b1;
  else
    Yb7l85 <= Oas675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nd7l85 <= 1'b1;
  else
    Nd7l85 <= Cbs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cf7l85 <= 1'b1;
  else
    Cf7l85 <= Cfv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rg7l85 <= 1'b1;
  else
    Rg7l85 <= Ghv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gi7l85 <= 1'b1;
  else
    Gi7l85 <= Uhv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vj7l85 <= 1'b1;
  else
    Vj7l85 <= Wiv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kl7l85 <= 1'b0;
  else
    Kl7l85 <= Xkx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zm7l85 <= 1'b0;
  else
    Zm7l85 <= Oyw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qo7l85 <= 1'b0;
  else
    Qo7l85 <= Hyw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hq7l85 <= 1'b0;
  else
    Hq7l85 <= Txw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yr7l85 <= 1'b0;
  else
    Yr7l85 <= Mxw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pt7l85 <= 1'b0;
  else
    Pt7l85 <= Fxw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gv7l85 <= 1'b0;
  else
    Gv7l85 <= Ypw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xw7l85 <= 1'b0;
  else
    Xw7l85 <= Rpw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Oy7l85 <= 1'b0;
  else
    Oy7l85 <= Dpw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    F08l85 <= 1'b0;
  else
    F08l85 <= Wow675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    W18l85 <= 1'b0;
  else
    W18l85 <= Pow675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    N38l85 <= 1'b0;
  else
    N38l85 <= F0q675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    E58l85 <= 1'b1;
  else
    E58l85 <= Nwu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    T68l85 <= 1'b1;
  else
    T68l85 <= Ryu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I88l85 <= 1'b1;
  else
    I88l85 <= Fzu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    X98l85 <= 1'b0;
  else
    X98l85 <= Paw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ib8l85 <= 1'b1;
  else
    Ib8l85 <= Xxr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xc8l85 <= 1'b0;
  else
    Xc8l85 <= Qxr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ke8l85 <= 1'b0;
  else
    Ke8l85 <= Jxr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xf8l85 <= 1'b0;
  else
    Xf8l85 <= Cxr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kh8l85 <= 1'b1;
  else
    Kh8l85 <= S1w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yi8l85 <= 1'b0;
  else
    Yi8l85 <= Pux675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jk8l85 <= 1'b1;
  else
    Jk8l85 <= Xmv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xl8l85 <= 1'b1;
  else
    Xl8l85 <= Ppv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ln8l85 <= 1'b1;
  else
    Ln8l85 <= Wux675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zo8l85 <= 1'b1;
  else
    Zo8l85 <= Twx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nq8l85 <= 1'b0;
  else
    Nq8l85 <= F3y675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Es8l85 <= 1'b0;
  else
    Es8l85 <= Amp675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vt8l85 <= 1'b1;
  else
    Vt8l85 <= Pdt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kv8l85 <= 1'b1;
  else
    Kv8l85 <= Tft675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zw8l85 <= 1'b1;
  else
    Zw8l85 <= Hgt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Oy8l85 <= 1'b1;
  else
    Oy8l85 <= Jht675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    D09l85 <= 1'b0;
  else
    D09l85 <= Mbq675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    V19l85 <= 1'b1;
  else
    V19l85 <= Zcs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    J39l85 <= 1'b1;
  else
    J39l85 <= Dfs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    X49l85 <= 1'b1;
  else
    X49l85 <= Rfs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    L69l85 <= 1'b1;
  else
    L69l85 <= Tgs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Z79l85 <= 1'b0;
  else
    Z79l85 <= Qyp675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Q99l85 <= 1'b1;
  else
    Q99l85 <= Zsx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Eb9l85 <= 1'b1;
  else
    Eb9l85 <= Kox675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sc9l85 <= 1'b1;
  else
    Sc9l85 <= Bux675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ge9l85 <= 1'b1;
  else
    Ge9l85 <= X9u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Uf9l85 <= 1'b1;
  else
    Uf9l85 <= Bcu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ih9l85 <= 1'b1;
  else
    Ih9l85 <= Pcu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wi9l85 <= 1'b1;
  else
    Wi9l85 <= Rdu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kk9l85 <= 1'b1;
  else
    Kk9l85 <= Q6x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bm9l85 <= 1'b1;
  else
    Bm9l85 <= L0x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sn9l85 <= 1'b1;
  else
    Sn9l85 <= O5x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ip9l85 <= 1'b1;
  else
    Ip9l85 <= H5x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yq9l85 <= 1'b1;
  else
    Yq9l85 <= Eit675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ns9l85 <= 1'b1;
  else
    Ns9l85 <= Ikt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cu9l85 <= 1'b1;
  else
    Cu9l85 <= Wkt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rv9l85 <= 1'b1;
  else
    Rv9l85 <= Ylt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gx9l85 <= 1'b1;
  else
    Gx9l85 <= E7x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xy9l85 <= 1'b1;
  else
    Xy9l85 <= Z0x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    O0al85 <= 1'b1;
  else
    O0al85 <= Eqs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    B2al85 <= 1'b1;
  else
    B2al85 <= Pls675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    P3al85 <= 1'b1;
  else
    P3al85 <= I9x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    F5al85 <= 1'b1;
  else
    F5al85 <= D3x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    V6al85 <= 1'b1;
  else
    V6al85 <= Qzw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    M8al85 <= 1'b1;
  else
    M8al85 <= Qnu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Aaal85 <= 1'b1;
  else
    Aaal85 <= Upu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Obal85 <= 1'b1;
  else
    Obal85 <= Iqu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cdal85 <= 1'b1;
  else
    Cdal85 <= Kru675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qeal85 <= 1'b0;
  else
    Qeal85 <= Ayw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hgal85 <= 1'b0;
  else
    Hgal85 <= Kpw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yhal85 <= 1'b0;
  else
    Yhal85 <= Ngw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mjal85 <= 1'b1;
  else
    Mjal85 <= Qrx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Alal85 <= 1'b1;
  else
    Alal85 <= Vwr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Omal85 <= 1'b1;
  else
    Omal85 <= Bju675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Coal85 <= 1'b1;
  else
    Coal85 <= Flu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qpal85 <= 1'b1;
  else
    Qpal85 <= Tlu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Eral85 <= 1'b1;
  else
    Eral85 <= Vmu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ssal85 <= 1'b1;
  else
    Ssal85 <= C6x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jual85 <= 1'b1;
  else
    Jual85 <= Xzw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Awal85 <= 1'b1;
  else
    Awal85 <= Gav675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pxal85 <= 1'b1;
  else
    Pxal85 <= Kcv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ezal85 <= 1'b1;
  else
    Ezal85 <= Ycv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    T0bl85 <= 1'b1;
  else
    T0bl85 <= Aev675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I2bl85 <= 1'b0;
  else
    I2bl85 <= Mwq675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    A4bl85 <= 1'b0;
  else
    A4bl85 <= Qew675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    L5bl85 <= 1'b0;
  else
    L5bl85 <= L8w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    D7bl85 <= 1'b0;
  else
    D7bl85 <= K3q675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    V8bl85 <= 1'b1;
  else
    V8bl85 <= R5v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kabl85 <= 1'b1;
  else
    Kabl85 <= V7v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zbbl85 <= 1'b1;
  else
    Zbbl85 <= J8v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Odbl85 <= 1'b1;
  else
    Odbl85 <= L9v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dfbl85 <= 1'b0;
  else
    Dfbl85 <= Gtq675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vgbl85 <= 1'b1;
  else
    Vgbl85 <= Irt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kibl85 <= 1'b1;
  else
    Kibl85 <= Mtt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zjbl85 <= 1'b1;
  else
    Zjbl85 <= Aut675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Olbl85 <= 1'b1;
  else
    Olbl85 <= Xvt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dnbl85 <= 1'b1;
  else
    Dnbl85 <= Byt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sobl85 <= 1'b1;
  else
    Sobl85 <= Pyt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hqbl85 <= 1'b1;
  else
    Hqbl85 <= M0u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wrbl85 <= 1'b1;
  else
    Wrbl85 <= Q2u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ltbl85 <= 1'b1;
  else
    Ltbl85 <= E3u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Avbl85 <= 1'b1;
  else
    Avbl85 <= C1v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pwbl85 <= 1'b1;
  else
    Pwbl85 <= G3v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Eybl85 <= 1'b1;
  else
    Eybl85 <= U3v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tzbl85 <= 1'b1;
  else
    Tzbl85 <= W4v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I1cl85 <= 1'b0;
  else
    I1cl85 <= Qrq675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    A3cl85 <= 1'b1;
  else
    A3cl85 <= Tmt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    P4cl85 <= 1'b1;
  else
    P4cl85 <= Xot675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    E6cl85 <= 1'b1;
  else
    E6cl85 <= Lpt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    T7cl85 <= 1'b1;
  else
    T7cl85 <= Nqt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I9cl85 <= 1'b0;
  else
    I9cl85 <= Seq675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Abcl85 <= 1'b1;
  else
    Abcl85 <= Xrx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Occl85 <= 1'b1;
  else
    Occl85 <= Esx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cecl85 <= 1'b0;
  else
    Cecl85 <= Y2y675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qfcl85 <= 1'b0;
  else
    Qfcl85 <= Owr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dhcl85 <= 1'b0;
  else
    Dhcl85 <= Utx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qicl85 <= 1'b1;
  else
    Qicl85 <= Gtx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bkcl85 <= 1'b0;
  else
    Bkcl85 <= A6w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nlcl85 <= 1'b1;
  else
    Nlcl85 <= Jrx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bncl85 <= 1'b1;
  else
    Bncl85 <= Crx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pocl85 <= 1'b1;
  else
    Pocl85 <= Vqx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dqcl85 <= 1'b1;
  else
    Dqcl85 <= Oqx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rrcl85 <= 1'b1;
  else
    Rrcl85 <= Hqx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gtcl85 <= 1'b1;
  else
    Gtcl85 <= Aqx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vucl85 <= 1'b1;
  else
    Vucl85 <= Tpx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kwcl85 <= 1'b1;
  else
    Kwcl85 <= Mpx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zxcl85 <= 1'b1;
  else
    Zxcl85 <= Z1w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nzcl85 <= 1'b1;
  else
    Nzcl85 <= Hwr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Z0dl85 <= 1'b1;
  else
    Z0dl85 <= Awr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    L2dl85 <= 1'b0;
  else
    L2dl85 <= W1y675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    B4dl85 <= 1'b0;
  else
    B4dl85 <= Iaw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    N5dl85 <= 1'b0;
  else
    N5dl85 <= Gjp675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Z6dl85 <= 1'b0;
  else
    Z6dl85 <= Mcw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    L8dl85 <= 1'b0;
  else
    L8dl85 <= Ihw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cadl85 <= 1'b1;
  else
    Cadl85 <= I3w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ubdl85 <= 1'b0;
  else
    Ubdl85 <= Tvr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Iddl85 <= 1'b1;
  else
    Iddl85 <= Mvr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xedl85 <= 1'b1;
  else
    Xedl85 <= Fvr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lgdl85 <= 1'b1;
  else
    Lgdl85 <= Yur675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zhdl85 <= 1'b1;
  else
    Zhdl85 <= Rur675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Njdl85 <= 1'b1;
  else
    Njdl85 <= Kur675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bldl85 <= 1'b1;
  else
    Bldl85 <= Dur675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pmdl85 <= 1'b1;
  else
    Pmdl85 <= Wtr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dodl85 <= 1'b1;
  else
    Dodl85 <= Ptr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rpdl85 <= 1'b1;
  else
    Rpdl85 <= Itr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Frdl85 <= 1'b1;
  else
    Frdl85 <= Btr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tsdl85 <= 1'b1;
  else
    Tsdl85 <= Usr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hudl85 <= 1'b1;
  else
    Hudl85 <= Nsr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wvdl85 <= 1'b1;
  else
    Wvdl85 <= Gsr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lxdl85 <= 1'b1;
  else
    Lxdl85 <= Zrr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Azdl85 <= 1'b1;
  else
    Azdl85 <= Srr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    P0el85 <= 1'b1;
  else
    P0el85 <= Lrr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    E2el85 <= 1'b1;
  else
    E2el85 <= Err675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    T3el85 <= 1'b1;
  else
    T3el85 <= Szx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I5el85 <= 1'b1;
  else
    I5el85 <= Xqr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    W6el85 <= 1'b0;
  else
    W6el85 <= Fwx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    K8el85 <= 1'b0;
  else
    K8el85 <= Qqr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Y9el85 <= 1'b0;
  else
    Y9el85 <= Whw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nbel85 <= 1'b0;
  else
    Nbel85 <= Czw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Edel85 <= 1'b0;
  else
    Edel85 <= Mqw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Veel85 <= 1'b0;
  else
    Veel85 <= Vyw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mgel85 <= 1'b0;
  else
    Mgel85 <= Fqw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Diel85 <= 1'b0;
  else
    Diel85 <= Baw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pjel85 <= 1'b0;
  else
    Pjel85 <= Jqr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Clel85 <= 1'b1;
  else
    Clel85 <= Cqr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nmel85 <= 1'b0;
  else
    Nmel85 <= Y4w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Znel85 <= 1'b1;
  else
    Znel85 <= Vpr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kpel85 <= 1'b1;
  else
    Kpel85 <= Opr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vqel85 <= 1'b1;
  else
    Vqel85 <= Hpr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gsel85 <= 1'b1;
  else
    Gsel85 <= Apr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rtel85 <= 1'b1;
  else
    Rtel85 <= Tor675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cvel85 <= 1'b1;
  else
    Cvel85 <= Mor675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nwel85 <= 1'b1;
  else
    Nwel85 <= For675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yxel85 <= 1'b1;
  else
    Yxel85 <= Ynr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kzel85 <= 1'b1;
  else
    Kzel85 <= Rnr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    W0fl85 <= 1'b1;
  else
    W0fl85 <= Knr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I2fl85 <= 1'b1;
  else
    I2fl85 <= Dnr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    U3fl85 <= 1'b1;
  else
    U3fl85 <= Wmr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    G5fl85 <= 1'b1;
  else
    G5fl85 <= Pmr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    S6fl85 <= 1'b1;
  else
    S6fl85 <= Imr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    E8fl85 <= 1'b1;
  else
    E8fl85 <= Bmr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Q9fl85 <= 1'b1;
  else
    Q9fl85 <= Ulr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cbfl85 <= 1'b1;
  else
    Cbfl85 <= Nlr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ocfl85 <= 1'b1;
  else
    Ocfl85 <= Glr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Aefl85 <= 1'b1;
  else
    Aefl85 <= Zkr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mffl85 <= 1'b1;
  else
    Mffl85 <= Skr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ygfl85 <= 1'b1;
  else
    Ygfl85 <= Lkr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kifl85 <= 1'b1;
  else
    Kifl85 <= Ekr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wjfl85 <= 1'b1;
  else
    Wjfl85 <= Xjr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ilfl85 <= 1'b1;
  else
    Ilfl85 <= Dox675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wmfl85 <= 1'b1;
  else
    Wmfl85 <= Wnx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kofl85 <= 1'b1;
  else
    Kofl85 <= Pnx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ypfl85 <= 1'b1;
  else
    Ypfl85 <= Inx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mrfl85 <= 1'b1;
  else
    Mrfl85 <= Bnx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Atfl85 <= 1'b1;
  else
    Atfl85 <= Umx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Oufl85 <= 1'b1;
  else
    Oufl85 <= Nmx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cwfl85 <= 1'b1;
  else
    Cwfl85 <= Gmx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qxfl85 <= 1'b1;
  else
    Qxfl85 <= Zlx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fzfl85 <= 1'b1;
  else
    Fzfl85 <= Slx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    U0gl85 <= 1'b1;
  else
    U0gl85 <= Llx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    J2gl85 <= 1'b1;
  else
    J2gl85 <= Tkv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    U3gl85 <= 1'b1;
  else
    U3gl85 <= B3w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    M5gl85 <= 1'b1;
  else
    M5gl85 <= U2w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    E7gl85 <= 1'b1;
  else
    E7gl85 <= N2w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    W8gl85 <= 1'b1;
  else
    W8gl85 <= Qjr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kagl85 <= 1'b1;
  else
    Kagl85 <= Jjr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ybgl85 <= 1'b1;
  else
    Ybgl85 <= Cjr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mdgl85 <= 1'b1;
  else
    Mdgl85 <= Vir675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Afgl85 <= 1'b1;
  else
    Afgl85 <= Oir675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Oggl85 <= 1'b1;
  else
    Oggl85 <= Ipv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Digl85 <= 1'b1;
  else
    Digl85 <= Bpv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sjgl85 <= 1'b1;
  else
    Sjgl85 <= Uov675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Glgl85 <= 1'b1;
  else
    Glgl85 <= Nov675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Umgl85 <= 1'b1;
  else
    Umgl85 <= Gov675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Iogl85 <= 1'b1;
  else
    Iogl85 <= Nhv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xpgl85 <= 1'b1;
  else
    Xpgl85 <= Rcv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mrgl85 <= 1'b1;
  else
    Mrgl85 <= C8v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Btgl85 <= 1'b1;
  else
    Btgl85 <= N3v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qugl85 <= 1'b1;
  else
    Qugl85 <= Yyu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fwgl85 <= 1'b1;
  else
    Fwgl85 <= Quu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Uxgl85 <= 1'b1;
  else
    Uxgl85 <= Bqu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Izgl85 <= 1'b1;
  else
    Izgl85 <= Mlu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    W0hl85 <= 1'b1;
  else
    W0hl85 <= Xgu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    K2hl85 <= 1'b1;
  else
    K2hl85 <= Icu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Y3hl85 <= 1'b1;
  else
    Y3hl85 <= X2u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    N5hl85 <= 1'b1;
  else
    N5hl85 <= Iyt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    C7hl85 <= 1'b1;
  else
    C7hl85 <= Ttt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    R8hl85 <= 1'b1;
  else
    R8hl85 <= Ept675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gahl85 <= 1'b1;
  else
    Gahl85 <= Pkt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vbhl85 <= 1'b1;
  else
    Vbhl85 <= Agt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kdhl85 <= 1'b1;
  else
    Kdhl85 <= Lbt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zehl85 <= 1'b1;
  else
    Zehl85 <= Oos675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nghl85 <= 1'b1;
  else
    Nghl85 <= Kfs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bihl85 <= 1'b1;
  else
    Bihl85 <= Vas675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qjhl85 <= 1'b1;
  else
    Qjhl85 <= Qmv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Flhl85 <= 1'b1;
  else
    Flhl85 <= Jmv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Umhl85 <= 1'b1;
  else
    Umhl85 <= Cmv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Iohl85 <= 1'b1;
  else
    Iohl85 <= Vlv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wphl85 <= 1'b1;
  else
    Wphl85 <= Olv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Krhl85 <= 1'b1;
  else
    Krhl85 <= Zgv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zshl85 <= 1'b1;
  else
    Zshl85 <= Dcv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ouhl85 <= 1'b1;
  else
    Ouhl85 <= O7v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dwhl85 <= 1'b1;
  else
    Dwhl85 <= Z2v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sxhl85 <= 1'b1;
  else
    Sxhl85 <= Kyu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hzhl85 <= 1'b1;
  else
    Hzhl85 <= Cuu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    W0il85 <= 1'b1;
  else
    W0il85 <= Npu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    K2il85 <= 1'b1;
  else
    K2il85 <= Yku675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Y3il85 <= 1'b1;
  else
    Y3il85 <= Jgu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    M5il85 <= 1'b1;
  else
    M5il85 <= Ubu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    A7il85 <= 1'b1;
  else
    A7il85 <= J2u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    P8il85 <= 1'b1;
  else
    P8il85 <= Uxt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Eail85 <= 1'b1;
  else
    Eail85 <= Ftt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tbil85 <= 1'b1;
  else
    Tbil85 <= Qot675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Idil85 <= 1'b1;
  else
    Idil85 <= Bkt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xeil85 <= 1'b1;
  else
    Xeil85 <= Mft675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mgil85 <= 1'b1;
  else
    Mgil85 <= Xat675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Biil85 <= 1'b1;
  else
    Biil85 <= Aos675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pjil85 <= 1'b1;
  else
    Pjil85 <= Wes675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dlil85 <= 1'b1;
  else
    Dlil85 <= Has675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Smil85 <= 1'b1;
  else
    Smil85 <= Rjv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Goil85 <= 1'b1;
  else
    Goil85 <= Kjv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vpil85 <= 1'b1;
  else
    Vpil85 <= Djv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kril85 <= 1'b1;
  else
    Kril85 <= Piv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zsil85 <= 1'b1;
  else
    Zsil85 <= Tdv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ouil85 <= 1'b1;
  else
    Ouil85 <= E9v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dwil85 <= 1'b1;
  else
    Dwil85 <= P4v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sxil85 <= 1'b1;
  else
    Sxil85 <= Svu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hzil85 <= 1'b1;
  else
    Hzil85 <= Dru675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    V0jl85 <= 1'b1;
  else
    V0jl85 <= Omu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    J2jl85 <= 1'b1;
  else
    J2jl85 <= Zhu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    X3jl85 <= 1'b1;
  else
    X3jl85 <= Kdu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    L5jl85 <= 1'b1;
  else
    L5jl85 <= Gqt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    A7jl85 <= 1'b1;
  else
    A7jl85 <= Rlt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    P8jl85 <= 1'b1;
  else
    P8jl85 <= Cht675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Eajl85 <= 1'b1;
  else
    Eajl85 <= Nct675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tbjl85 <= 1'b1;
  else
    Tbjl85 <= Qps675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hdjl85 <= 1'b1;
  else
    Hdjl85 <= Mgs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vejl85 <= 1'b1;
  else
    Vejl85 <= Mkv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jgjl85 <= 1'b1;
  else
    Jgjl85 <= Fkv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yhjl85 <= 1'b1;
  else
    Yhjl85 <= Yjv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Njjl85 <= 1'b1;
  else
    Njjl85 <= Asv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cljl85 <= 1'b1;
  else
    Cljl85 <= Trv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rmjl85 <= 1'b1;
  else
    Rmjl85 <= Mrv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fojl85 <= 1'b1;
  else
    Fojl85 <= Frv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tpjl85 <= 1'b1;
  else
    Tpjl85 <= Yqv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hrjl85 <= 1'b1;
  else
    Hrjl85 <= Biv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wsjl85 <= 1'b1;
  else
    Wsjl85 <= Fdv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lujl85 <= 1'b1;
  else
    Lujl85 <= Q8v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Awjl85 <= 1'b1;
  else
    Awjl85 <= B4v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pxjl85 <= 1'b1;
  else
    Pxjl85 <= Evu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ezjl85 <= 1'b1;
  else
    Ezjl85 <= Pqu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    S0kl85 <= 1'b1;
  else
    S0kl85 <= Amu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    G2kl85 <= 1'b1;
  else
    G2kl85 <= Lhu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    U3kl85 <= 1'b1;
  else
    U3kl85 <= Wcu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I5kl85 <= 1'b1;
  else
    I5kl85 <= Spt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    X6kl85 <= 1'b1;
  else
    X6kl85 <= Dlt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    M8kl85 <= 1'b1;
  else
    M8kl85 <= Ogt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bakl85 <= 1'b1;
  else
    Bakl85 <= Zbt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qbkl85 <= 1'b1;
  else
    Qbkl85 <= Cps675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Edkl85 <= 1'b1;
  else
    Edkl85 <= Yfs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sekl85 <= 1'b1;
  else
    Sekl85 <= Jtv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hgkl85 <= 1'b1;
  else
    Hgkl85 <= Ctv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Whkl85 <= 1'b1;
  else
    Whkl85 <= Vsv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kjkl85 <= 1'b1;
  else
    Kjkl85 <= Osv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ykkl85 <= 1'b1;
  else
    Ykkl85 <= Hsv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mmkl85 <= 1'b1;
  else
    Mmkl85 <= Iiv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bokl85 <= 1'b1;
  else
    Bokl85 <= Mdv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qpkl85 <= 1'b1;
  else
    Qpkl85 <= X8v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Frkl85 <= 1'b1;
  else
    Frkl85 <= I4v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Uskl85 <= 1'b1;
  else
    Uskl85 <= Lvu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jukl85 <= 1'b1;
  else
    Jukl85 <= Wqu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xvkl85 <= 1'b1;
  else
    Xvkl85 <= Hmu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lxkl85 <= 1'b1;
  else
    Lxkl85 <= Shu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zykl85 <= 1'b1;
  else
    Zykl85 <= Ddu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    N0ll85 <= 1'b1;
  else
    N0ll85 <= Zpt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    C2ll85 <= 1'b1;
  else
    C2ll85 <= Klt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    R3ll85 <= 1'b1;
  else
    R3ll85 <= Vgt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    G5ll85 <= 1'b1;
  else
    G5ll85 <= Gct675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    V6ll85 <= 1'b1;
  else
    V6ll85 <= Jps675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    J8ll85 <= 1'b1;
  else
    J8ll85 <= Fgs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    X9ll85 <= 1'b1;
  else
    X9ll85 <= Suv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mbll85 <= 1'b1;
  else
    Mbll85 <= Luv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bdll85 <= 1'b1;
  else
    Bdll85 <= Euv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pell85 <= 1'b1;
  else
    Pell85 <= Xtv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dgll85 <= 1'b1;
  else
    Dgll85 <= Qtv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rhll85 <= 1'b1;
  else
    Rhll85 <= Sgv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gjll85 <= 1'b1;
  else
    Gjll85 <= Wbv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vkll85 <= 1'b1;
  else
    Vkll85 <= H7v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kmll85 <= 1'b1;
  else
    Kmll85 <= S2v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Znll85 <= 1'b1;
  else
    Znll85 <= Dyu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Opll85 <= 1'b1;
  else
    Opll85 <= Vtu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Drll85 <= 1'b1;
  else
    Drll85 <= Gpu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rsll85 <= 1'b1;
  else
    Rsll85 <= Rku675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Full85 <= 1'b1;
  else
    Full85 <= Cgu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tvll85 <= 1'b1;
  else
    Tvll85 <= Nbu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hxll85 <= 1'b1;
  else
    Hxll85 <= C2u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wyll85 <= 1'b1;
  else
    Wyll85 <= Nxt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    L0ml85 <= 1'b1;
  else
    L0ml85 <= Yst675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    A2ml85 <= 1'b1;
  else
    A2ml85 <= Jot675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    P3ml85 <= 1'b1;
  else
    P3ml85 <= Ujt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    E5ml85 <= 1'b1;
  else
    E5ml85 <= Fft675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    T6ml85 <= 1'b1;
  else
    T6ml85 <= Qat675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I8ml85 <= 1'b1;
  else
    I8ml85 <= Tns675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    W9ml85 <= 1'b1;
  else
    W9ml85 <= Pes675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kbml85 <= 1'b1;
  else
    Kbml85 <= Aas675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zcml85 <= 1'b1;
  else
    Zcml85 <= Bwv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Oeml85 <= 1'b1;
  else
    Oeml85 <= Uvv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dgml85 <= 1'b1;
  else
    Dgml85 <= Nvv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rhml85 <= 1'b1;
  else
    Rhml85 <= Gvv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fjml85 <= 1'b1;
  else
    Fjml85 <= Zuv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tkml85 <= 1'b1;
  else
    Tkml85 <= Lgv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Imml85 <= 1'b1;
  else
    Imml85 <= Pbv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xnml85 <= 1'b1;
  else
    Xnml85 <= A7v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mpml85 <= 1'b1;
  else
    Mpml85 <= L2v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Brml85 <= 1'b1;
  else
    Brml85 <= Wxu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qsml85 <= 1'b1;
  else
    Qsml85 <= Otu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fuml85 <= 1'b1;
  else
    Fuml85 <= Zou675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tvml85 <= 1'b1;
  else
    Tvml85 <= Kku675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hxml85 <= 1'b1;
  else
    Hxml85 <= Vfu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vyml85 <= 1'b1;
  else
    Vyml85 <= Gbu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    J0nl85 <= 1'b1;
  else
    J0nl85 <= V1u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Y1nl85 <= 1'b1;
  else
    Y1nl85 <= Gxt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    N3nl85 <= 1'b1;
  else
    N3nl85 <= Rst675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    C5nl85 <= 1'b1;
  else
    C5nl85 <= Cot675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    R6nl85 <= 1'b1;
  else
    R6nl85 <= Njt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    G8nl85 <= 1'b1;
  else
    G8nl85 <= Yet675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    V9nl85 <= 1'b1;
  else
    V9nl85 <= Jat675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kbnl85 <= 1'b1;
  else
    Kbnl85 <= Mns675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ycnl85 <= 1'b1;
  else
    Ycnl85 <= Ies675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Menl85 <= 1'b1;
  else
    Menl85 <= T9s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bgnl85 <= 1'b1;
  else
    Bgnl85 <= Kxv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qhnl85 <= 1'b1;
  else
    Qhnl85 <= Dxv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fjnl85 <= 1'b1;
  else
    Fjnl85 <= Wwv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tknl85 <= 1'b1;
  else
    Tknl85 <= Pwv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hmnl85 <= 1'b1;
  else
    Hmnl85 <= Iwv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vnnl85 <= 1'b1;
  else
    Vnnl85 <= Egv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kpnl85 <= 1'b1;
  else
    Kpnl85 <= Ibv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zqnl85 <= 1'b1;
  else
    Zqnl85 <= T6v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Osnl85 <= 1'b1;
  else
    Osnl85 <= E2v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dunl85 <= 1'b1;
  else
    Dunl85 <= Pxu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Svnl85 <= 1'b1;
  else
    Svnl85 <= Htu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hxnl85 <= 1'b1;
  else
    Hxnl85 <= Sou675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vynl85 <= 1'b1;
  else
    Vynl85 <= Dku675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    J0ol85 <= 1'b1;
  else
    J0ol85 <= Ofu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    X1ol85 <= 1'b1;
  else
    X1ol85 <= Zau675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    L3ol85 <= 1'b1;
  else
    L3ol85 <= O1u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    A5ol85 <= 1'b1;
  else
    A5ol85 <= Zwt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    P6ol85 <= 1'b1;
  else
    P6ol85 <= Kst675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    E8ol85 <= 1'b1;
  else
    E8ol85 <= Vnt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    T9ol85 <= 1'b1;
  else
    T9ol85 <= Gjt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ibol85 <= 1'b1;
  else
    Ibol85 <= Ret675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xcol85 <= 1'b1;
  else
    Xcol85 <= Cat675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Meol85 <= 1'b1;
  else
    Meol85 <= Fns675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Agol85 <= 1'b1;
  else
    Agol85 <= Bes675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ohol85 <= 1'b1;
  else
    Ohol85 <= M9s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Djol85 <= 1'b1;
  else
    Djol85 <= Tyv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Skol85 <= 1'b1;
  else
    Skol85 <= Myv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hmol85 <= 1'b1;
  else
    Hmol85 <= Fyv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vnol85 <= 1'b1;
  else
    Vnol85 <= Yxv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jpol85 <= 1'b1;
  else
    Jpol85 <= Rxv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xqol85 <= 1'b1;
  else
    Xqol85 <= Xfv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Msol85 <= 1'b1;
  else
    Msol85 <= Bbv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Buol85 <= 1'b1;
  else
    Buol85 <= M6v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qvol85 <= 1'b1;
  else
    Qvol85 <= X1v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fxol85 <= 1'b1;
  else
    Fxol85 <= Ixu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Uyol85 <= 1'b1;
  else
    Uyol85 <= Atu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    J0pl85 <= 1'b1;
  else
    J0pl85 <= Lou675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    X1pl85 <= 1'b1;
  else
    X1pl85 <= Wju675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    L3pl85 <= 1'b1;
  else
    L3pl85 <= Hfu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Z4pl85 <= 1'b1;
  else
    Z4pl85 <= Sau675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    N6pl85 <= 1'b1;
  else
    N6pl85 <= H1u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    C8pl85 <= 1'b1;
  else
    C8pl85 <= Swt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    R9pl85 <= 1'b1;
  else
    R9pl85 <= Dst675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gbpl85 <= 1'b1;
  else
    Gbpl85 <= Ont675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vcpl85 <= 1'b1;
  else
    Vcpl85 <= Zit675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kepl85 <= 1'b1;
  else
    Kepl85 <= Ket675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zfpl85 <= 1'b1;
  else
    Zfpl85 <= V9t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ohpl85 <= 1'b1;
  else
    Ohpl85 <= Yms675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cjpl85 <= 1'b1;
  else
    Cjpl85 <= Uds675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qkpl85 <= 1'b1;
  else
    Qkpl85 <= F9s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fmpl85 <= 1'b1;
  else
    Fmpl85 <= C0w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Unpl85 <= 1'b1;
  else
    Unpl85 <= Vzv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jppl85 <= 1'b1;
  else
    Jppl85 <= Ozv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xqpl85 <= 1'b1;
  else
    Xqpl85 <= Hzv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lspl85 <= 1'b1;
  else
    Lspl85 <= Azv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ztpl85 <= 1'b1;
  else
    Ztpl85 <= Qfv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ovpl85 <= 1'b1;
  else
    Ovpl85 <= Uav675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dxpl85 <= 1'b1;
  else
    Dxpl85 <= F6v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sypl85 <= 1'b1;
  else
    Sypl85 <= Q1v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    H0ql85 <= 1'b1;
  else
    H0ql85 <= Bxu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    W1ql85 <= 1'b1;
  else
    W1ql85 <= Tsu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    L3ql85 <= 1'b1;
  else
    L3ql85 <= Eou675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Z4ql85 <= 1'b1;
  else
    Z4ql85 <= Pju675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    N6ql85 <= 1'b1;
  else
    N6ql85 <= Afu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    B8ql85 <= 1'b1;
  else
    B8ql85 <= Lau675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    P9ql85 <= 1'b1;
  else
    P9ql85 <= A1u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ebql85 <= 1'b1;
  else
    Ebql85 <= Lwt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tcql85 <= 1'b1;
  else
    Tcql85 <= Wrt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ieql85 <= 1'b1;
  else
    Ieql85 <= Hnt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xfql85 <= 1'b1;
  else
    Xfql85 <= Sit675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mhql85 <= 1'b1;
  else
    Mhql85 <= Det675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bjql85 <= 1'b1;
  else
    Bjql85 <= O9t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qkql85 <= 1'b1;
  else
    Qkql85 <= Rms675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Emql85 <= 1'b1;
  else
    Emql85 <= Nds675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Snql85 <= 1'b1;
  else
    Snql85 <= Y8s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hpql85 <= 1'b1;
  else
    Hpql85 <= L1w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wqql85 <= 1'b1;
  else
    Wqql85 <= E1w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lsql85 <= 1'b1;
  else
    Lsql85 <= X0w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ztql85 <= 1'b1;
  else
    Ztql85 <= Q0w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nvql85 <= 1'b1;
  else
    Nvql85 <= J0w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bxql85 <= 1'b1;
  else
    Bxql85 <= Jfv675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qyql85 <= 1'b1;
  else
    Qyql85 <= Nav675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    F0rl85 <= 1'b1;
  else
    F0rl85 <= Y5v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    U1rl85 <= 1'b1;
  else
    U1rl85 <= J1v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    J3rl85 <= 1'b1;
  else
    J3rl85 <= Uwu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Y4rl85 <= 1'b1;
  else
    Y4rl85 <= Msu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    N6rl85 <= 1'b1;
  else
    N6rl85 <= Xnu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    B8rl85 <= 1'b1;
  else
    B8rl85 <= Iju675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    P9rl85 <= 1'b1;
  else
    P9rl85 <= Teu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dbrl85 <= 1'b1;
  else
    Dbrl85 <= Eau675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rcrl85 <= 1'b1;
  else
    Rcrl85 <= T0u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gerl85 <= 1'b1;
  else
    Gerl85 <= Ewt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vfrl85 <= 1'b1;
  else
    Vfrl85 <= Prt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Khrl85 <= 1'b1;
  else
    Khrl85 <= Ant675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zirl85 <= 1'b1;
  else
    Zirl85 <= Lit675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Okrl85 <= 1'b1;
  else
    Okrl85 <= Wdt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dmrl85 <= 1'b1;
  else
    Dmrl85 <= H9t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Snrl85 <= 1'b1;
  else
    Snrl85 <= Kms675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gprl85 <= 1'b1;
  else
    Gprl85 <= Gds675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Uqrl85 <= 1'b1;
  else
    Uqrl85 <= R8s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jsrl85 <= 1'b1;
  else
    Jsrl85 <= Vev675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ytrl85 <= 1'b1;
  else
    Ytrl85 <= Z9v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nvrl85 <= 1'b1;
  else
    Nvrl85 <= K5v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cxrl85 <= 1'b1;
  else
    Cxrl85 <= V0v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ryrl85 <= 1'b1;
  else
    Ryrl85 <= Gwu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    G0sl85 <= 1'b1;
  else
    G0sl85 <= Yru675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    V1sl85 <= 1'b1;
  else
    V1sl85 <= Jnu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    J3sl85 <= 1'b1;
  else
    J3sl85 <= Uiu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    X4sl85 <= 1'b1;
  else
    X4sl85 <= Feu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    L6sl85 <= 1'b1;
  else
    L6sl85 <= Q9u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Z7sl85 <= 1'b1;
  else
    Z7sl85 <= Ydu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    N9sl85 <= 1'b1;
  else
    N9sl85 <= F0u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cbsl85 <= 1'b1;
  else
    Cbsl85 <= Qvt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rcsl85 <= 1'b1;
  else
    Rcsl85 <= Brt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gesl85 <= 1'b1;
  else
    Gesl85 <= Mmt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vfsl85 <= 1'b1;
  else
    Vfsl85 <= Xht675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Khsl85 <= 1'b1;
  else
    Khsl85 <= Idt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zisl85 <= 1'b1;
  else
    Zisl85 <= T8t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Oksl85 <= 1'b1;
  else
    Oksl85 <= Wls675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cmsl85 <= 1'b1;
  else
    Cmsl85 <= W3w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qnsl85 <= 1'b1;
  else
    Qnsl85 <= Hhs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Epsl85 <= 1'b1;
  else
    Epsl85 <= Ohs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sqsl85 <= 1'b1;
  else
    Sqsl85 <= Vhs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gssl85 <= 1'b1;
  else
    Gssl85 <= Cis675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Utsl85 <= 1'b1;
  else
    Utsl85 <= Jis675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ivsl85 <= 1'b1;
  else
    Ivsl85 <= Qis675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wwsl85 <= 1'b1;
  else
    Wwsl85 <= Xis675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kysl85 <= 1'b1;
  else
    Kysl85 <= Ejs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yzsl85 <= 1'b1;
  else
    Yzsl85 <= Ljs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    M1tl85 <= 1'b1;
  else
    M1tl85 <= Sjs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    A3tl85 <= 1'b1;
  else
    A3tl85 <= Zjs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    O4tl85 <= 1'b1;
  else
    O4tl85 <= Gks675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    C6tl85 <= 1'b1;
  else
    C6tl85 <= Nks675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Q7tl85 <= 1'b1;
  else
    Q7tl85 <= Uks675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    E9tl85 <= 1'b1;
  else
    E9tl85 <= Bls675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Satl85 <= 1'b1;
  else
    Satl85 <= Ils675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gctl85 <= 1'b1;
  else
    Gctl85 <= Scs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Udtl85 <= 1'b1;
  else
    Udtl85 <= D8s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jftl85 <= 1'b0;
  else
    Jftl85 <= Mwx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zgtl85 <= 1'b1;
  else
    Zgtl85 <= P3w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nitl85 <= 1'b1;
  else
    Nitl85 <= Hir675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bktl85 <= 1'b1;
  else
    Bktl85 <= Air675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nltl85 <= 1'b1;
  else
    Nltl85 <= O3s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cntl85 <= 1'b1;
  else
    Cntl85 <= C4s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rotl85 <= 1'b1;
  else
    Rotl85 <= J4s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gqtl85 <= 1'b1;
  else
    Gqtl85 <= Q4s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vrtl85 <= 1'b1;
  else
    Vrtl85 <= X4s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kttl85 <= 1'b1;
  else
    Kttl85 <= E5s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zutl85 <= 1'b1;
  else
    Zutl85 <= L5s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Owtl85 <= 1'b1;
  else
    Owtl85 <= S5s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dytl85 <= 1'b1;
  else
    Dytl85 <= Z5s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sztl85 <= 1'b1;
  else
    Sztl85 <= G6s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    H1ul85 <= 1'b1;
  else
    H1ul85 <= U6s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    W2ul85 <= 1'b1;
  else
    W2ul85 <= B7s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    L4ul85 <= 1'b1;
  else
    L4ul85 <= I7s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    A6ul85 <= 1'b1;
  else
    A6ul85 <= P7s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    P7ul85 <= 1'b0;
  else
    P7ul85 <= Zfw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    F9ul85 <= 1'b0;
  else
    F9ul85 <= Sfw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vaul85 <= 1'b1;
  else
    Vaul85 <= Cnu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jcul85 <= 1'b1;
  else
    Jcul85 <= Rru675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xdul85 <= 1'b1;
  else
    Xdul85 <= Hxx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lful85 <= 1'b1;
  else
    Lful85 <= Ahs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zgul85 <= 1'b0;
  else
    Zgul85 <= P1y675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Piul85 <= 1'b0;
  else
    Piul85 <= Vcx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ekul85 <= 1'b0;
  else
    Ekul85 <= Jdx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tlul85 <= 1'b0;
  else
    Tlul85 <= Qdx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Inul85 <= 1'b0;
  else
    Inul85 <= Xdx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xoul85 <= 1'b0;
  else
    Xoul85 <= Eex675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mqul85 <= 1'b0;
  else
    Mqul85 <= Lex675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bsul85 <= 1'b0;
  else
    Bsul85 <= Sex675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qtul85 <= 1'b0;
  else
    Qtul85 <= Zex675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fvul85 <= 1'b0;
  else
    Fvul85 <= Gfx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vwul85 <= 1'b0;
  else
    Vwul85 <= Igx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lyul85 <= 1'b0;
  else
    Lyul85 <= Pgx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    B0vl85 <= 1'b0;
  else
    B0vl85 <= Wgx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    R1vl85 <= 1'b0;
  else
    R1vl85 <= Dhx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    H3vl85 <= 1'b0;
  else
    H3vl85 <= Khx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    X4vl85 <= 1'b0;
  else
    X4vl85 <= Rhx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    N6vl85 <= 1'b0;
  else
    N6vl85 <= Yhx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    D8vl85 <= 1'b0;
  else
    D8vl85 <= Fix675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    T9vl85 <= 1'b0;
  else
    T9vl85 <= Mix675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jbvl85 <= 1'b0;
  else
    Jbvl85 <= Tix675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zcvl85 <= 1'b0;
  else
    Zcvl85 <= Ajx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pevl85 <= 1'b0;
  else
    Pevl85 <= Hjx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fgvl85 <= 1'b0;
  else
    Fgvl85 <= Ojx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vhvl85 <= 1'b0;
  else
    Vhvl85 <= Vjx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ljvl85 <= 1'b0;
  else
    Ljvl85 <= Ckx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Blvl85 <= 1'b0;
  else
    Blvl85 <= Jkx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rmvl85 <= 1'b0;
  else
    Rmvl85 <= Qkx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hovl85 <= 1'b0;
  else
    Hovl85 <= U0y675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wpvl85 <= 1'b0;
  else
    Wpvl85 <= B1y675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mrvl85 <= 1'b0;
  else
    Mrvl85 <= Bhw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Atvl85 <= 1'b0;
  else
    Atvl85 <= Ugw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ouvl85 <= 1'b0;
  else
    Ouvl85 <= Phw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cwvl85 <= 1'b0;
  else
    Cwvl85 <= Cdx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rxvl85 <= 1'b0;
  else
    Rxvl85 <= Clw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Izvl85 <= 1'b0;
  else
    Izvl85 <= Emw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Y0wl85 <= 1'b0;
  else
    Y0wl85 <= Xlw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    O2wl85 <= 1'b0;
  else
    O2wl85 <= Qlw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    F4wl85 <= 1'b0;
  else
    F4wl85 <= Jlw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    W5wl85 <= 1'b0;
  else
    W5wl85 <= Vkw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    N7wl85 <= 1'b0;
  else
    N7wl85 <= Okw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    E9wl85 <= 1'b0;
  else
    E9wl85 <= Hkw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vawl85 <= 1'b0;
  else
    Vawl85 <= Yiw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lcwl85 <= 1'b0;
  else
    Lcwl85 <= Akw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bewl85 <= 1'b0;
  else
    Bewl85 <= Tjw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rfwl85 <= 1'b0;
  else
    Rfwl85 <= Mjw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hhwl85 <= 1'b0;
  else
    Hhwl85 <= Fjw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xiwl85 <= 1'b0;
  else
    Xiwl85 <= Riw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nkwl85 <= 1'b0;
  else
    Nkwl85 <= Kiw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dmwl85 <= 1'b0;
  else
    Dmwl85 <= Diw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tnwl85 <= 1'b0;
  else
    Tnwl85 <= Stw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kpwl85 <= 1'b0;
  else
    Kpwl85 <= Uuw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Brwl85 <= 1'b0;
  else
    Brwl85 <= Nuw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sswl85 <= 1'b0;
  else
    Sswl85 <= Guw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Juwl85 <= 1'b0;
  else
    Juwl85 <= Ztw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Awwl85 <= 1'b0;
  else
    Awwl85 <= Ltw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rxwl85 <= 1'b0;
  else
    Rxwl85 <= Etw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Izwl85 <= 1'b0;
  else
    Izwl85 <= Xsw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Z0xl85 <= 1'b0;
  else
    Z0xl85 <= Orw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Q2xl85 <= 1'b0;
  else
    Q2xl85 <= Qsw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    H4xl85 <= 1'b0;
  else
    H4xl85 <= Jsw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Y5xl85 <= 1'b0;
  else
    Y5xl85 <= Csw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    P7xl85 <= 1'b0;
  else
    P7xl85 <= Vrw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    G9xl85 <= 1'b0;
  else
    G9xl85 <= Hrw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xaxl85 <= 1'b0;
  else
    Xaxl85 <= Arw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ocxl85 <= 1'b0;
  else
    Ocxl85 <= Tqw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fexl85 <= 1'b0;
  else
    Fexl85 <= Gnw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wfxl85 <= 1'b0;
  else
    Wfxl85 <= Iow675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nhxl85 <= 1'b0;
  else
    Nhxl85 <= Bow675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ejxl85 <= 1'b0;
  else
    Ejxl85 <= Unw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vkxl85 <= 1'b0;
  else
    Vkxl85 <= Nnw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mmxl85 <= 1'b0;
  else
    Mmxl85 <= Zmw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Doxl85 <= 1'b0;
  else
    Doxl85 <= Smw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Upxl85 <= 1'b0;
  else
    Upxl85 <= Lmw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lrxl85 <= 1'b0;
  else
    Lrxl85 <= D4w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dtxl85 <= 1'b0;
  else
    Dtxl85 <= K4w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vuxl85 <= 1'b0;
  else
    Vuxl85 <= R4w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nwxl85 <= 1'b0;
  else
    Nwxl85 <= Cdq675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fyxl85 <= 1'b0;
  else
    Fyxl85 <= M5w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wzxl85 <= 1'b0;
  else
    Wzxl85 <= Pnp675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    N1yl85 <= 1'b0;
  else
    N1yl85 <= T5w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    E3yl85 <= 1'b0;
  else
    E3yl85 <= Epp675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    V4yl85 <= 1'b0;
  else
    V4yl85 <= H6w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    N6yl85 <= 1'b0;
  else
    N6yl85 <= V6w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    F8yl85 <= 1'b0;
  else
    F8yl85 <= C7w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    X9yl85 <= 1'b0;
  else
    X9yl85 <= J7w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pbyl85 <= 1'b0;
  else
    Pbyl85 <= Q7w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gdyl85 <= 1'b0;
  else
    Gdyl85 <= E8w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yeyl85 <= 1'b0;
  else
    Yeyl85 <= G9w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qgyl85 <= 1'b0;
  else
    Qgyl85 <= N9w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Iiyl85 <= 1'b0;
  else
    Iiyl85 <= Waw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zjyl85 <= 1'b0;
  else
    Zjyl85 <= Tqp675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qlyl85 <= 1'b0;
  else
    Qlyl85 <= Dbw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hnyl85 <= 1'b0;
  else
    Hnyl85 <= Isp675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yoyl85 <= 1'b0;
  else
    Yoyl85 <= Kbw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pqyl85 <= 1'b0;
  else
    Pqyl85 <= Xtp675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gsyl85 <= 1'b0;
  else
    Gsyl85 <= Rbw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xtyl85 <= 1'b0;
  else
    Xtyl85 <= Mvp675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ovyl85 <= 1'b0;
  else
    Ovyl85 <= Ybw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fxyl85 <= 1'b0;
  else
    Fxyl85 <= Bxp675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wyyl85 <= 1'b0;
  else
    Wyyl85 <= Tcw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    O0zl85 <= 1'b0;
  else
    O0zl85 <= Adw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    G2zl85 <= 1'b0;
  else
    G2zl85 <= Ojq675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Y3zl85 <= 1'b0;
  else
    Y3zl85 <= Hdw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Q5zl85 <= 1'b0;
  else
    Q5zl85 <= Elq675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I7zl85 <= 1'b0;
  else
    I7zl85 <= Odw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    A9zl85 <= 1'b0;
  else
    A9zl85 <= Umq675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sazl85 <= 1'b0;
  else
    Sazl85 <= Cew675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kczl85 <= 1'b0;
  else
    Kczl85 <= Jew675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cezl85 <= 1'b0;
  else
    Cezl85 <= Igq675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ufzl85 <= 1'b0;
  else
    Ufzl85 <= Xew675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mhzl85 <= 1'b0;
  else
    Mhzl85 <= Efw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ejzl85 <= 1'b0;
  else
    Ejzl85 <= Wvw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vkzl85 <= 1'b0;
  else
    Vkzl85 <= Yww675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mmzl85 <= 1'b0;
  else
    Mmzl85 <= Rww675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dozl85 <= 1'b0;
  else
    Dozl85 <= Kww675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Upzl85 <= 1'b0;
  else
    Upzl85 <= Dww675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lrzl85 <= 1'b0;
  else
    Lrzl85 <= Pvw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ctzl85 <= 1'b0;
  else
    Ctzl85 <= Ivw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tuzl85 <= 1'b0;
  else
    Tuzl85 <= Bvw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kwzl85 <= 1'b0;
  else
    Kwzl85 <= Ocx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ayzl85 <= 1'b0;
  else
    Ayzl85 <= Hcx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rzzl85 <= 1'b0;
  else
    Rzzl85 <= Acx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I10m85 <= 1'b0;
  else
    I10m85 <= F5w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    W20m85 <= 1'b0;
  else
    W20m85 <= Lfw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    K40m85 <= 1'b1;
  else
    K40m85 <= V5x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    B60m85 <= 1'b1;
  else
    B60m85 <= T3y675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    S70m85 <= 1'b1;
  else
    S70m85 <= Tbx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I90m85 <= 1'b1;
  else
    I90m85 <= Mbx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ya0m85 <= 1'b1;
  else
    Ya0m85 <= Fbx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Oc0m85 <= 1'b1;
  else
    Oc0m85 <= A5x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ee0m85 <= 1'b1;
  else
    Ee0m85 <= Thr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pf0m85 <= 1'b1;
  else
    Pf0m85 <= Yax675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fh0m85 <= 1'b1;
  else
    Fh0m85 <= T4x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vi0m85 <= 1'b1;
  else
    Vi0m85 <= Rax675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lk0m85 <= 1'b1;
  else
    Lk0m85 <= M4x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bm0m85 <= 1'b1;
  else
    Bm0m85 <= Kax675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rn0m85 <= 1'b1;
  else
    Rn0m85 <= F4x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hp0m85 <= 1'b1;
  else
    Hp0m85 <= Dax675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xq0m85 <= 1'b1;
  else
    Xq0m85 <= Y3x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ns0m85 <= 1'b1;
  else
    Ns0m85 <= W9x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Du0m85 <= 1'b1;
  else
    Du0m85 <= R3x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tv0m85 <= 1'b1;
  else
    Tv0m85 <= P9x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jx0m85 <= 1'b1;
  else
    Jx0m85 <= K3x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zy0m85 <= 1'b1;
  else
    Zy0m85 <= B9x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Q01m85 <= 1'b1;
  else
    Q01m85 <= W2x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    H21m85 <= 1'b1;
  else
    H21m85 <= Z7x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Y31m85 <= 1'b1;
  else
    Y31m85 <= U1x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    P51m85 <= 1'b1;
  else
    P51m85 <= S7x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    G71m85 <= 1'b1;
  else
    G71m85 <= N1x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    X81m85 <= 1'b1;
  else
    X81m85 <= L7x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Oa1m85 <= 1'b1;
  else
    Oa1m85 <= G1x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fc1m85 <= 1'b1;
  else
    Fc1m85 <= X6x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wd1m85 <= 1'b1;
  else
    Wd1m85 <= S0x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nf1m85 <= 1'b1;
  else
    Nf1m85 <= J6x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Eh1m85 <= 1'b1;
  else
    Eh1m85 <= E0x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vi1m85 <= 1'b1;
  else
    Vi1m85 <= Tus675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kk1m85 <= 1'b1;
  else
    Kk1m85 <= Lqs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zl1m85 <= 1'b1;
  else
    Zl1m85 <= Sqs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    On1m85 <= 1'b1;
  else
    On1m85 <= Zqs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dp1m85 <= 1'b1;
  else
    Dp1m85 <= Grs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sq1m85 <= 1'b1;
  else
    Sq1m85 <= Nrs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hs1m85 <= 1'b1;
  else
    Hs1m85 <= Urs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wt1m85 <= 1'b1;
  else
    Wt1m85 <= Bss675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lv1m85 <= 1'b1;
  else
    Lv1m85 <= Iss675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ax1m85 <= 1'b1;
  else
    Ax1m85 <= Pss675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Py1m85 <= 1'b1;
  else
    Py1m85 <= Wss675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    E02m85 <= 1'b1;
  else
    E02m85 <= Dts675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    T12m85 <= 1'b1;
  else
    T12m85 <= Kts675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I32m85 <= 1'b1;
  else
    I32m85 <= Mhr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    U42m85 <= 1'b1;
  else
    U42m85 <= Rts675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    J62m85 <= 1'b1;
  else
    J62m85 <= Yts675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Y72m85 <= 1'b1;
  else
    Y72m85 <= Fus675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    M92m85 <= 1'b1;
  else
    M92m85 <= Mus675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ab2m85 <= 1'b1;
  else
    Ab2m85 <= Izs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pc2m85 <= 1'b1;
  else
    Pc2m85 <= Avs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ee2m85 <= 1'b1;
  else
    Ee2m85 <= Hvs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tf2m85 <= 1'b1;
  else
    Tf2m85 <= Ovs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ih2m85 <= 1'b1;
  else
    Ih2m85 <= Vvs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xi2m85 <= 1'b1;
  else
    Xi2m85 <= Cws675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mk2m85 <= 1'b1;
  else
    Mk2m85 <= Jws675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bm2m85 <= 1'b1;
  else
    Bm2m85 <= Qws675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qn2m85 <= 1'b1;
  else
    Qn2m85 <= Xws675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fp2m85 <= 1'b1;
  else
    Fp2m85 <= Exs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Uq2m85 <= 1'b1;
  else
    Uq2m85 <= Lxs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Js2m85 <= 1'b1;
  else
    Js2m85 <= Sxs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yt2m85 <= 1'b1;
  else
    Yt2m85 <= Zxs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nv2m85 <= 1'b1;
  else
    Nv2m85 <= Fhr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zw2m85 <= 1'b1;
  else
    Zw2m85 <= Gys675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Oy2m85 <= 1'b1;
  else
    Oy2m85 <= Nys675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    D03m85 <= 1'b1;
  else
    D03m85 <= Uys675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    R13m85 <= 1'b1;
  else
    R13m85 <= Bzs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    F33m85 <= 1'b0;
  else
    F33m85 <= Nfx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    V43m85 <= 1'b1;
  else
    V43m85 <= U8x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    M63m85 <= 1'b1;
  else
    M63m85 <= P2x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    D83m85 <= 1'b1;
  else
    D83m85 <= X3t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    S93m85 <= 1'b1;
  else
    S93m85 <= Pzs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hb3m85 <= 1'b1;
  else
    Hb3m85 <= Wzs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wc3m85 <= 1'b1;
  else
    Wc3m85 <= D0t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Le3m85 <= 1'b1;
  else
    Le3m85 <= K0t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ag3m85 <= 1'b1;
  else
    Ag3m85 <= R0t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ph3m85 <= 1'b1;
  else
    Ph3m85 <= Y0t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ej3m85 <= 1'b1;
  else
    Ej3m85 <= F1t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tk3m85 <= 1'b1;
  else
    Tk3m85 <= M1t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Im3m85 <= 1'b1;
  else
    Im3m85 <= T1t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xn3m85 <= 1'b1;
  else
    Xn3m85 <= A2t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mp3m85 <= 1'b1;
  else
    Mp3m85 <= H2t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Br3m85 <= 1'b1;
  else
    Br3m85 <= O2t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qs3m85 <= 1'b1;
  else
    Qs3m85 <= Ygr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cu3m85 <= 1'b1;
  else
    Cu3m85 <= V2t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rv3m85 <= 1'b1;
  else
    Rv3m85 <= C3t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gx3m85 <= 1'b1;
  else
    Gx3m85 <= J3t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vy3m85 <= 1'b1;
  else
    Vy3m85 <= Q3t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    K04m85 <= 1'b0;
  else
    K04m85 <= Ufx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    A24m85 <= 1'b1;
  else
    A24m85 <= N8x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    R34m85 <= 1'b1;
  else
    R34m85 <= I2x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I54m85 <= 1'b0;
  else
    I54m85 <= S8w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    A74m85 <= 1'b0;
  else
    A74m85 <= A5q675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    S84m85 <= 1'b1;
  else
    S84m85 <= M8t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ha4m85 <= 1'b1;
  else
    Ha4m85 <= E4t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wb4m85 <= 1'b1;
  else
    Wb4m85 <= L4t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ld4m85 <= 1'b1;
  else
    Ld4m85 <= S4t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Af4m85 <= 1'b1;
  else
    Af4m85 <= Z4t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pg4m85 <= 1'b1;
  else
    Pg4m85 <= G5t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ei4m85 <= 1'b1;
  else
    Ei4m85 <= N5t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tj4m85 <= 1'b1;
  else
    Tj4m85 <= U5t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Il4m85 <= 1'b1;
  else
    Il4m85 <= B6t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xm4m85 <= 1'b1;
  else
    Xm4m85 <= I6t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mo4m85 <= 1'b1;
  else
    Mo4m85 <= P6t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bq4m85 <= 1'b1;
  else
    Bq4m85 <= W6t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qr4m85 <= 1'b1;
  else
    Qr4m85 <= D7t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ft4m85 <= 1'b1;
  else
    Ft4m85 <= K7t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Uu4m85 <= 1'b1;
  else
    Uu4m85 <= R7t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jw4m85 <= 1'b1;
  else
    Jw4m85 <= Y7t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yx4m85 <= 1'b1;
  else
    Yx4m85 <= F8t675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nz4m85 <= 1'b0;
  else
    Nz4m85 <= Bgx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    D15m85 <= 1'b1;
  else
    D15m85 <= G8x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    U25m85 <= 1'b1;
  else
    U25m85 <= B2x675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    L45m85 <= 1'b0;
  else
    L45m85 <= Z8w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    D65m85 <= 1'b0;
  else
    D65m85 <= Q6q675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    V75m85 <= 1'b1;
  else
    V75m85 <= Bdt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    K95m85 <= 1'b1;
  else
    K95m85 <= Qht675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Za5m85 <= 1'b1;
  else
    Za5m85 <= Fmt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Oc5m85 <= 1'b1;
  else
    Oc5m85 <= Uqt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    De5m85 <= 1'b1;
  else
    De5m85 <= N0y675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sf5m85 <= 1'b1;
  else
    Sf5m85 <= D5v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hh5m85 <= 1'b1;
  else
    Hh5m85 <= S9v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wi5m85 <= 1'b1;
  else
    Wi5m85 <= Cyx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lk5m85 <= 1'b1;
  else
    Lk5m85 <= Qyx675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Am5m85 <= 1'b1;
  else
    Am5m85 <= A3s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pn5m85 <= 1'b1;
  else
    Pn5m85 <= Rgr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bp5m85 <= 1'b1;
  else
    Bp5m85 <= U4u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qq5m85 <= 1'b1;
  else
    Qq5m85 <= B5u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fs5m85 <= 1'b1;
  else
    Fs5m85 <= I5u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ut5m85 <= 1'b1;
  else
    Ut5m85 <= P5u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jv5m85 <= 1'b1;
  else
    Jv5m85 <= W5u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yw5m85 <= 1'b1;
  else
    Yw5m85 <= D6u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ny5m85 <= 1'b1;
  else
    Ny5m85 <= K6u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    C06m85 <= 1'b1;
  else
    C06m85 <= R6u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    R16m85 <= 1'b1;
  else
    R16m85 <= Y6u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    G36m85 <= 1'b1;
  else
    G36m85 <= F7u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    V46m85 <= 1'b1;
  else
    V46m85 <= M7u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    K66m85 <= 1'b1;
  else
    K66m85 <= T7u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Z76m85 <= 1'b1;
  else
    Z76m85 <= A8u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    O96m85 <= 1'b1;
  else
    O96m85 <= H8u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Db6m85 <= 1'b1;
  else
    Db6m85 <= O8u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sc6m85 <= 1'b1;
  else
    Sc6m85 <= V8u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    He6m85 <= 1'b1;
  else
    He6m85 <= C9u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wf6m85 <= 1'b1;
  else
    Wf6m85 <= L3u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lh6m85 <= 1'b1;
  else
    Lh6m85 <= S3u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Aj6m85 <= 1'b1;
  else
    Aj6m85 <= Z3u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pk6m85 <= 1'b1;
  else
    Pk6m85 <= G4u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Em6m85 <= 1'b1;
  else
    Em6m85 <= N4u675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tn6m85 <= 1'b1;
  else
    Tn6m85 <= Wyt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ip6m85 <= 1'b1;
  else
    Ip6m85 <= Dzt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xq6m85 <= 1'b1;
  else
    Xq6m85 <= Kzt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ms6m85 <= 1'b1;
  else
    Ms6m85 <= Rzt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bu6m85 <= 1'b1;
  else
    Bu6m85 <= Yzt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qv6m85 <= 1'b1;
  else
    Qv6m85 <= Hut675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fx6m85 <= 1'b1;
  else
    Fx6m85 <= Out675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Uy6m85 <= 1'b1;
  else
    Uy6m85 <= Vut675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    J07m85 <= 1'b1;
  else
    J07m85 <= Cvt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Y17m85 <= 1'b1;
  else
    Y17m85 <= Jvt675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    N37m85 <= 1'b1;
  else
    N37m85 <= Jzw675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    E57m85 <= 1'b0;
  else
    E57m85 <= X7w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    V67m85 <= 1'b0;
  else
    V67m85 <= O6w675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    N87m85 <= 1'b1;
  else
    N87m85 <= Mzu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ca7m85 <= 1'b1;
  else
    Ca7m85 <= Tzu675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rb7m85 <= 1'b1;
  else
    Rb7m85 <= A0v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gd7m85 <= 1'b1;
  else
    Gd7m85 <= H0v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ve7m85 <= 1'b1;
  else
    Ve7m85 <= O0v675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kg7m85 <= 1'b1;
  else
    Kg7m85 <= Jbs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zh7m85 <= 1'b1;
  else
    Zh7m85 <= Qbs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Oj7m85 <= 1'b1;
  else
    Oj7m85 <= Xbs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dl7m85 <= 1'b1;
  else
    Dl7m85 <= Ecs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sm7m85 <= 1'b1;
  else
    Sm7m85 <= Lcs675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ho7m85 <= 1'b0;
  else
    Ho7m85 <= Kgr675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xp7m85 <= 1'b1;
  else
    Xp7m85 <= W7s675;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mr7m85 <= 1'b0;
  else
    Mr7m85 <= Dgr675;

endmodule

//------------------------------------------------------------------------------
// EOF
//------------------------------------------------------------------------------

